module invader_ROM (
	
	input clk,
	input resetN,
	input [31:0] adress, // for future purpose
	output [15:0] dout,
	output [17:0] depth,
	output [31:0] repeats

);



/* invader killing sound*/
 // stroe the value
bit [0:3376][15:0] invader_ROM ={ // need to be 0 to 102 so first 2 bytes be on the left 
16'h0000, 16'h0000, 16'h0001, 16'hFFFE,
 16'h0002, 16'hFFFE, 16'h0002, 16'h0000,
 16'hFFFF, 16'h0000, 16'h0000, 16'h0000,
 16'h0002, 16'hFFFD, 16'h0002, 16'hFFFE,
 16'h0003, 16'hFFFD, 16'h0002, 16'hFFFE,
 16'h0001, 16'h0001, 16'hFFFF, 16'h0000,
 16'h0001, 16'hFFFE, 16'h0001, 16'h0001,
 16'hFFFF, 16'h0000, 16'h0001, 16'hFFFE,
 16'h0003, 16'hFFFD, 16'h0002, 16'hFFFF,
 16'h0001, 16'hFFFF, 16'h0000, 16'h0001,
 16'hFFFF, 16'h0001, 16'hFFFF, 16'h0000,
 16'h0001, 16'hFFFF, 16'h0001, 16'hFFFF,
 16'h0001, 16'hFFFE, 16'h0004, 16'hFFFB,
 16'h0004, 16'hFFFE, 16'h0000, 16'h0002,
 16'hFFFD, 16'h0003, 16'hFFFD, 16'h0003,
 16'hFFFD, 16'h0003, 16'hFFFD, 16'h0002,
 16'hFFFF, 16'h0001, 16'hFFFE, 16'h0003,
 16'hFFFC, 16'h0005, 16'hFFFC, 16'h0002,
 16'hFFFF, 16'h0001, 16'hFFFF, 16'h0001,
 16'hFFFF, 16'h0001, 16'h0000, 16'hFFFF,
 16'h0001, 16'hFFFF, 16'h0001, 16'h0000,
 16'h0000, 16'h0000, 16'h0000, 16'hFFFF,
 16'h0002, 16'hFFFD, 16'h0004, 16'hFFFC,
 16'h0003, 16'hFFFD, 16'h0003, 16'hFFFD,
 16'h1004, 16'h23FA, 16'h1109, 16'hEEF4,
 16'hDF10, 16'hDAEC, 16'hE417, 16'hE9E6,
 16'hFE1E, 16'h05DE, 16'hEC28, 16'hECD1,
 16'hFB36, 16'h1FC3, 16'h1E44, 16'hF5B5,
 16'hE553, 16'h0FA5, 16'h3D62, 16'hED98,
 16'hCF6D, 16'h198F, 16'h4A76, 16'hF483,
 16'h9083, 16'hDF78, 16'h508C, 16'h3A72,
 16'hC18F, 16'hE36F, 16'h4093, 16'h2E6C,
 16'hDD93, 16'h8000, 16'hEA8D, 16'h7C77,
 16'h0984, 16'h9082, 16'h0C77, 16'h7190,
 16'hE769, 16'h809E, 16'h065A, 16'h7EB0,
 16'h0645, 16'h83C6, 16'hEE2E, 16'h65DE,
 16'hF616, 16'h80F6, 16'h1500, 16'h7F08,
 16'hD8EF, 16'h861A, 16'h1FDE, 16'h7F2A,
 16'hEDCE, 16'h8038, 16'hBBC5, 16'h313C,
 16'h7EC5, 16'hD137, 16'h9ACF, 16'h4F29,
 16'h29E3, 16'hAB0E, 16'hBD03, 16'h47E9,
 16'h332E, 16'h96B8, 16'hE865, 16'h747C,
 16'hF0A4, 16'h8A3C, 16'hE6E4, 16'h50FB,
 16'h5A26, 16'hA5BB, 16'hCA63, 16'h6B81,
 16'hF398, 16'h9B52, 16'hBAC1, 16'h2B31,
 16'h7FFF, 16'hD925, 16'h81D9, 16'h0F2E,
 16'h7FFF, 16'h084D, 16'h8B9B, 16'hBC80,
 16'h2C60, 16'h7AC4, 16'hD515, 16'h8000,
 16'h2CBD, 16'h7370, 16'hAE62, 16'hAECB,
 16'h4F0A, 16'h3E20, 16'hC9B9, 16'h806B,
 16'h0C75, 16'h7FA6, 16'h1243, 16'h90CE,
 16'hC026, 16'h3FE2, 16'h561B, 16'h9EE2,
 16'hD325, 16'h60D0, 16'h223D, 16'hCEB4,
 16'h8000, 16'h0091, 16'h7E82, 16'hFC6B,
 16'h8000, 16'h154C, 16'h7EC0, 16'hE637,
 16'h8000, 16'h0A2B, 16'h78D6, 16'h292C,
 16'hBECE, 16'h803C, 16'h25B8, 16'h7F55,
 16'hBD9E, 16'h986F, 16'h4283, 16'h658A,
 16'hA06B, 16'hCE9F, 16'h5F5A, 16'h23AA,
 16'hC555, 16'h80A8, 16'h1060, 16'h7F92,
 16'hE382, 16'h8065, 16'h20B9, 16'h7F24,
 16'hDC04, 16'h8001, 16'h2361, 16'h7E6D,
 16'hDFC6, 16'h8000, 16'h072B, 16'h74A4,
 16'h408A, 16'hCB4B, 16'h81DC, 16'hFB03,
 16'h7FFF, 16'hFFCF, 16'h8240, 16'hD5B9,
 16'h4848, 16'h5FBF, 16'hE132, 16'h8001,
 16'hFC03, 16'h7D1D, 16'h1FBE, 16'hA96A,
 16'hB66B, 16'h53C3, 16'h330E, 16'h9420,
 16'hE3B5, 16'h5573, 16'h4869, 16'hB0B6,
 16'hA731, 16'h45E1, 16'h5615, 16'hCAED,
 16'h801A, 16'h02D5, 16'h7F46, 16'h0596,
 16'h8697, 16'hE734, 16'h5C08, 16'h31B5,
 16'h9395, 16'hE71C, 16'h7D36, 16'hE576,
 16'h86DE, 16'hE6D0, 16'h677F, 16'h4836,
 16'hB110, 16'hAEAF, 16'h3D8A, 16'h7248,
 16'hD0DA, 16'h8000, 16'h36F6, 16'h6F10,
 16'hABDC, 16'hAF46, 16'h4B8A, 16'h57B3,
 16'hD903, 16'h8000, 16'hEC48, 16'h7C28,
 16'h385E, 16'hA123, 16'hE456, 16'h7D36,
 16'hE03C, 16'h8053, 16'hF51E, 16'h506F,
 16'h7108, 16'hD67D, 16'h8001, 16'h0C74,
 16'h7B1F, 16'h0042, 16'h8000, 16'h10DF,
 16'h77E5, 16'hFE4A, 16'hA593, 16'h9883,
 16'h1C75, 16'h7FFF, 16'h0D8C, 16'h9458,
 16'hB6CE, 16'h3904, 16'h7A31, 16'hC293,
 16'h95B0, 16'h4808, 16'h5A44, 16'hDE6D,
 16'h8000, 16'h09CC, 16'h7C85, 16'hE22B,
 16'h8001, 16'h3390, 16'h7DB8, 16'hCD04,
 16'h853D, 16'h3386, 16'h7EB2, 16'hD01B,
 16'h8013, 16'h25C4, 16'h7F60, 16'hEB81,
 16'h8099, 16'hED53, 16'h7FBA, 16'hDB3F,
 16'h80C3, 16'hF940, 16'h64B7, 16'h5657,
 16'hB996, 16'h9782, 16'h3562, 16'h7BBD,
 16'hCB20, 16'h8005, 16'hF5D5, 16'h7F54,
 16'h0581, 16'h81AA, 16'h042B, 16'h56FF,
 16'h3ADB, 16'hC247, 16'h8000, 16'h247E,
 16'h7D6C, 16'hE0A6, 16'h8000, 16'h10BA,
 16'h7D46, 16'hFFB2, 16'hA05C, 16'hB190,
 16'h3F8A, 16'h7FFF, 16'hBFCF, 16'h9708,
 16'h4F24, 16'h49AC, 16'hB186, 16'h9F48,
 16'h50EA, 16'h46E6, 16'hAA46, 16'hC592,
 16'h3E92, 16'h7A4F, 16'hB9CA, 16'h8A23,
 16'h3EEA, 16'h5C10, 16'hD7EE, 16'h8001,
 16'h0CD6, 16'h7E40, 16'h01A4, 16'h9A7E,
 16'hD85A, 16'h50D3, 16'h49FC, 16'hB638,
 16'h9B94, 16'h3A9F, 16'h7A2E, 16'hDF03,
 16'h8000, 16'h115C, 16'h7D7D, 16'hD3A4,
 16'h8240, 16'h3FD6, 16'h7D1B, 16'hBDEC,
 16'h9115, 16'h4BE3, 16'h5A2C, 16'hABBD,
 16'hB561, 16'h557B, 16'h38AF, 16'hA421,
 16'hCD13, 16'h5DB5, 16'h2887, 16'h9B3B,
 16'hDF04, 16'h54BB, 16'h3D86, 16'hCA39,
 16'h8108, 16'h10BA, 16'h7FFF, 16'hEF49,
 16'h81EB, 16'h26E6, 16'h7FFF, 16'hD098,
 16'h8288, 16'hF35D, 16'h73B9, 16'h2135,
 16'h9BD7, 16'hE825, 16'h4CD8, 16'h512F,
 16'hD1C5, 16'h8003, 16'h07A1, 16'h7C76,
 16'h1B6E, 16'hA7B2, 16'hC02A, 16'h55FF,
 16'h25D5, 16'h8558, 16'h157A, 16'h63B6,
 16'h1B19, 16'hB519, 16'h80B3, 16'h3882,
 16'h7F49, 16'hC0EC, 16'h88DF, 16'h4555,
 16'h6779, 16'hB6B6, 16'hA11E, 16'h3E0C,
 16'h72CB, 16'hD15C, 16'h8005, 16'hF2A2,
 16'h6C40, 16'h53D9, 16'hA613, 16'hDBFC,
 16'h53FB, 16'h2108, 16'hB0F9, 16'h8402,
 16'h4308, 16'h5BE8, 16'hB92D, 16'hA0B8,
 16'h3E67, 16'h7FFF, 16'hC4AF, 16'h8928,
 16'h2703, 16'h7FD0, 16'hF95E, 16'h8075,
 16'hF4B7, 16'h6B1E, 16'hDC0B, 16'h86CF,
 16'h0253, 16'h6990, 16'h3C87, 16'h8F68,
 16'hFCA3, 16'h6459, 16'hF9A3, 16'hAD6A,
 16'h8F81, 16'h319C, 16'h7F40, 16'hE7EA,
 16'h8002, 16'h0E53, 16'h7E70, 16'hD7D1,
 16'h8000, 16'h1D5E, 16'h7C5B, 16'h04EC,
 16'h96CE, 16'hE676, 16'h5149, 16'h39F4,
 16'hBCD4, 16'h895D, 16'h207A, 16'h7FFF,
 16'hE73E, 16'h8BD5, 16'hDD20, 16'h36E2,
 16'h7B26, 16'hE6C8, 16'h8000, 16'hFC8C,
 16'h619A, 16'h1E3C, 16'hA8F3, 16'hD9DA,
 16'h535D, 16'h3769, 16'hB9D1, 16'hA4F6,
 16'h2D42, 16'h7FFF, 16'hF5A9, 16'h9027,
 16'hB105, 16'h27D5, 16'h7E4B, 16'hE29B,
 16'h8000, 16'h2B7D, 16'h708A, 16'hF174,
 16'h8D88, 16'hE17F, 16'h6D77, 16'hFF99,
 16'h9253, 16'h1FC2, 16'h7B26, 16'hDBF4,
 16'h8001, 16'h2326, 16'h79C1, 16'hFF56,
 16'h9394, 16'hE780, 16'h5271, 16'h2D9A,
 16'hBC5F, 16'h90A3, 16'h2C5F, 16'h7FFE,
 16'hD86E, 16'h8186, 16'h2189, 16'h6664,
 16'h27B2, 16'hB235, 16'h8CE7, 16'h3DFC,
 16'h6623, 16'hCEBC, 16'h8002, 16'h137C,
 16'h7EA3, 16'hFF40, 16'h9EDB, 16'hF80C,
 16'h5D0B, 16'h13E1, 16'hA430, 16'hD5C1,
 16'h634A, 16'hFEB0, 16'h9452, 16'h02B0,
 16'h5749, 16'h42C1, 16'hA632, 16'hC5DF,
 16'h4D0D, 16'h3209, 16'hC1DF, 16'h803B,
 16'h26A8, 16'h7F78, 16'hE668, 16'h85B7,
 16'h0A2A, 16'h57F2, 16'h2DF5, 16'hCA23,
 16'h8003, 16'h314C, 16'h7DA5, 16'hFB65,
 16'h8D97, 16'hE968, 16'h539D, 16'h2559,
 16'hC2B7, 16'h8133, 16'h31E8, 16'h7FF8,
 16'hC82C, 16'h96AB, 16'h4482, 16'h754D,
 16'hC0E7, 16'h8000, 16'h2F52, 16'h7E79,
 16'hD8BB, 16'h8000, 16'h281D, 16'h70B6,
 16'hF574, 16'hA567, 16'hAAB9, 16'h442B,
 16'h73EA, 16'hC107, 16'h8E03, 16'h28FA,
 16'h7FFF, 16'hE706, 16'h81EB, 16'h1329,
 16'h61BF, 16'h0C5D, 16'h9E85, 16'hD69C,
 16'h4441, 16'h44E3, 16'hBFF7, 16'h8000,
 16'h40AA, 16'h707B, 16'hC260, 16'h89C2,
 16'h3420, 16'h7EFB, 16'hD9EF, 16'h8022,
 16'h30CF, 16'h7A3D, 16'hBEBC, 16'h9847,
 16'h3EBA, 16'h6C40, 16'hD4C8, 16'h802F,
 16'h06DD, 16'h7713, 16'hE200, 16'h9CE9,
 16'h0630, 16'h5DB6, 16'h4565, 16'hB17F,
 16'hB49C, 16'h4749, 16'h51D3, 16'hB910,
 16'h940D, 16'h42D6, 16'h6747, 16'hB99D,
 16'h957D, 16'h2D6B, 16'h7FFF, 16'hE53D,
 16'h81D7, 16'h1C18, 16'h70F6, 16'hCDFE,
 16'h820C, 16'h11EE, 16'h5315, 16'h4BEA,
 16'hC912, 16'h8000, 16'h41FF, 16'h6810,
 16'hB9DD, 16'h9A38, 16'h3EB0, 16'h7D6B,
 16'hD678, 16'h8000, 16'h1636, 16'h6BED,
 16'h07EF, 16'hB236, 16'hA6A5, 16'h2D7F,
 16'h7F5E, 16'hDBC4, 16'h801D, 16'h10FE,
 16'h52EA, 16'h162B, 16'hBEC4, 16'h8749,
 16'h3CAE, 16'h7F56, 16'hBCAB, 16'h9150,
 16'h37B8, 16'h7F3D, 16'hF6D2, 16'h951B,
 16'hB3FC, 16'h35EA, 16'h7033, 16'hBEAF,
 16'h8070, 16'h3D70, 16'h75B0, 16'hD532,
 16'h84E9, 16'hFCFF, 16'h6616, 16'h27D7,
 16'hBF38, 16'hB5BD, 16'h444B, 16'h74B2,
 16'hB84B, 16'h8BBB, 16'h413B, 16'h71D5,
 16'hC217, 16'h8000, 16'h35E6, 16'h7A36,
 16'hF6AC, 16'hA974, 16'hA66A, 16'h3AB9,
 16'h7F25, 16'hC3FC, 16'h8001, 16'h3A38,
 16'h7EAD, 16'h036C, 16'hAC7F, 16'h9D93,
 16'h355E, 16'h7FAD, 16'hD24C, 16'h80B8,
 16'h1347, 16'h53B6, 16'h3A50, 16'hD1A8,
 16'h8000, 16'h3591, 16'h7E7E, 16'hD471,
 16'h88A0, 16'h1E4F, 16'h6FC1, 16'hDB31,
 16'h8ADD, 16'h3516, 16'h78F5, 16'hE301,
 16'h9308, 16'hF4F2, 16'h6512, 16'hEAED,
 16'hA111, 16'hF8F2, 16'h570A, 16'h4DFB,
 16'hA600, 16'hD707, 16'h54EF, 16'h191C,
 16'hAED8, 16'hAF35, 16'h52BF, 16'h314D,
 16'h9FA7, 16'hF764, 16'h6092, 16'h0078,
 16'h977F, 16'h1189, 16'h6B70, 16'hDB95,
 16'h9E68, 16'hF99A, 16'h4F65, 16'h579A,
 16'hBC68, 16'h8096, 16'h346E, 16'h7F8D,
 16'hD478, 16'h8282, 16'h2485, 16'h6476,
 16'hE28E, 16'h9C6D, 16'hDB99, 16'h5560,
 16'h41A7, 16'hA752, 16'hEBB3, 16'h534A,
 16'h23B9, 16'hC244, 16'h8000, 16'h3D40,
 16'h7EC4, 16'hED3A, 16'hA9C7, 16'hB538,
 16'h49C8, 16'h6339, 16'hBDC6, 16'h943C,
 16'h32C1, 16'h7F42, 16'hE2BC, 16'h9446,
 16'hE0B8, 16'h404A, 16'h5AB4, 16'hBB4E,
 16'h80B0, 16'h3E52, 16'h7EAC, 16'hD456,
 16'h96A8, 16'hD359, 16'h39A8, 16'h7F55,
 16'hBDAE, 16'h804F, 16'h3EB4, 16'h6C49,
 16'hC1BA, 16'h8041, 16'h40C6, 16'h7233,
 16'hBAD4, 16'h9C24, 16'h4FE3, 16'h5418,
 16'hB7ED, 16'h9E0E, 16'h34F5, 16'h7F09,
 16'hC0FA, 16'h8805, 16'h45F9, 16'h5D09,
 16'hADF3, 16'h9F14, 16'h4BE5, 16'h4B22,
 16'hA9D5, 16'hBF35, 16'h54C0, 16'h304D,
 16'hB4A6, 16'hB165, 16'h4191, 16'h7B79,
 16'hBB7E, 16'h868A, 16'h266F, 16'h7697,
 16'hDB65, 16'h939D, 16'h0463, 16'h479B,
 16'h5269, 16'hBC91, 16'h8002, 16'h2A7E,
 16'h7B8E, 16'hFE65, 16'h9FA8, 16'hE84B,
 16'h50C2, 16'h152F, 16'hA8E2, 16'hD10E,
 16'h4C00, 16'h3FF4, 16'hAA14, 16'hC9E8,
 16'h5A1A, 16'h1EE6, 16'hB118, 16'hC8EB,
 16'h4111, 16'h79F4, 16'hCE05, 16'h8003,
 16'h29F5, 16'h6B13, 16'hC2E7, 16'h8F1D,
 16'h30DF, 16'h7C23, 16'hD6DE, 16'h9F1F,
 16'hFDE8, 16'h430D, 16'h7301, 16'hC3ED,
 16'h8028, 16'h33C0, 16'h665C, 16'hBF87,
 16'h8897, 16'h1D49, 16'h72D7, 16'h010A,
 16'hA915, 16'hEBCD, 16'h404E, 16'h5D9A,
 16'hC17A, 16'h8002, 16'h2B93, 16'h6268,
 16'h1896, 16'hAD72, 16'hA780, 16'h4695,
 16'h5651, 16'hBDCD, 16'h8111, 16'h1715,
 16'h73C1, 16'h266D, 16'hA763, 16'hFBCE,
 16'h5E01, 16'hE92F, 16'hB5A3, 16'hAB89,
 16'h3D4F, 16'h7FD5, 16'hB80A, 16'h8F12,
 16'h2DD8, 16'h6C39, 16'h0CBC, 16'h9D48,
 16'hD9BA, 16'h433E, 16'h29D0, 16'hAF1D,
 16'h95FA, 16'h49EC, 16'h6F31, 16'hC5AF,
 16'h8673, 16'h0F69, 16'h6EBC, 16'h1120,
 16'hA203, 16'h1CDB, 16'h6E45, 16'hCE9D,
 16'hA97E, 16'hD56B, 16'h3EA8, 16'h7E49,
 16'hBBC2, 16'h8001, 16'h3FCE, 16'h6930,
 16'hF0D0, 16'hA733, 16'hABC6, 16'h4444,
 16'h78B0, 16'hB85E, 16'h8393, 16'h417C,
 16'h7F75, 16'hC599, 16'h9159, 16'h3EB5,
 16'h683F, 16'hD2CB, 16'h8D2C, 16'hEADB,
 16'h511F, 16'h3DE7, 16'hB614, 16'hA8EF,
 16'h510F, 16'h58F3, 16'hB40C, 16'h98F4,
 16'h4D0D, 16'h6EF1, 16'hB611, 16'h93ED,
 16'h4015, 16'h7AEA, 16'hF117, 16'h9CE8,
 16'hAB17, 16'h3DEC, 16'h7D11, 16'hB3F2,
 16'h800B, 16'h10F8, 16'h6B05, 16'h24FE,
 16'hA1FE, 16'h0505, 16'h5FFA, 16'hF407,
 16'hA0F8, 16'hDE07, 16'h53FB, 16'h2502,
 16'hA103, 16'hE2F7, 16'h6610, 16'hECE8,
 16'h9721, 16'h35D5, 16'h6935, 16'hEDC2,
 16'hA046, 16'hE9B4, 16'h5A4F, 16'h13B2,
 16'h9E4A, 16'hFFBD, 16'h6838, 16'hD5D7,
 16'h8F17, 16'h3F00, 16'h6FE4, 16'hE03B,
 16'hA9A2, 16'hC986, 16'h484E, 16'h7CE2,
 16'hABEB, 16'h8749, 16'h4E83, 16'h6FB1,
 16'hB31B, 16'h8219, 16'h1AB4, 16'h797B,
 16'hFF5B, 16'hABCA, 16'hE516, 16'h4105,
 16'h6FE5, 16'hAD2C, 16'h8000, 16'h333B,
 16'h5AC9, 16'h0F2D, 16'hA8E3, 16'h8907,
 16'h4614, 16'h7FFF, 16'hB657, 16'h8281,
 16'h26A9, 16'h5A2C, 16'h2D00, 16'hB2D3,
 16'h8E59, 16'h5A7C, 16'h49AF, 16'hA128,
 16'hC6FE, 16'h55DD, 16'h3847, 16'hAD98,
 16'hB286, 16'h6260, 16'h2FB6, 16'hA436,
 16'hD8DC, 16'h4913, 16'h79FD, 16'hC4F5,
 16'h8017, 16'h30DF, 16'h6328, 16'hB4D2,
 16'h9533, 16'h17C9, 16'h753B, 16'h14C1,
 16'hA743, 16'hDDB9, 16'h484B, 16'h79B1,
 16'hBB52, 16'h8000, 16'h0652, 16'h57AE,
 16'h1251, 16'h9AB0, 16'h104F, 16'h5FB4,
 16'hF947, 16'hACBE, 16'hAE3C, 16'h55CA,
 16'h7030, 16'h9ED7, 16'hC022, 16'h60E5,
 16'h1D14, 16'hA7F2, 16'hDB08, 16'h4CFF,
 16'h4DFA, 16'hAB0D, 16'h8FEC, 16'h541A,
 16'h7DE2, 16'hCB21, 16'h8000, 16'h2028,
 16'h6BD4, 16'hCE30, 16'hA4CC, 16'hF638,
 16'h56C5, 16'h573D, 16'hA2C1, 16'hC441,
 16'h50BB, 16'h444B, 16'hADAF, 16'h8257,
 16'h50A4, 16'h7160, 16'hBB9C, 16'h8169,
 16'h2D91, 16'h7975, 16'hCF86, 16'hA67F,
 16'h0A7D, 16'h5585, 16'h5C79, 16'hAB89,
 16'h8002, 16'h368A, 16'h7176, 16'h068A,
 16'h9377, 16'hE486, 16'h4C7E, 16'h217D,
 16'hB089, 16'h8572, 16'h5093, 16'h7F67,
 16'hAB9E, 16'hA25D, 16'h5EAA, 16'h5B50,
 16'hABB4, 16'h9549, 16'h3AB9, 16'h7F47,
 16'hBFB8, 16'h9948, 16'h07B9, 16'h6146,
 16'h27BC, 16'h8F42, 16'h05BF, 16'h4C41,
 16'h0ABE, 16'hA244, 16'hA3B9, 16'h524A,
 16'h5AB5, 16'hB24B, 16'h85B6, 16'h5847,
 16'h6CBC, 16'hA242, 16'hB9C1, 16'h513B,
 16'h5DCA, 16'hB530, 16'h8001, 16'h3C25,
 16'h65E0, 16'h0C1A, 16'hA3ED, 16'hC10C,
 16'h62FA, 16'h0E01, 16'hA903, 16'hD5F9,
 16'h5A0C, 16'h52EF, 16'h9D14, 16'hD1EB,
 16'h5A15, 16'h24EB, 16'hA515, 16'hB2E9,
 16'h4E1A, 16'h6EE4, 16'hA21D, 16'h82E2,
 16'h5C1F, 16'h55DF, 16'hA924, 16'hA0D9,
 16'h4B2A, 16'h7ED3, 16'hB631, 16'h83C9,
 16'h2C3F, 16'h67B8, 16'hE251, 16'h98A7,
 16'h1162, 16'h5394, 16'h0978, 16'h9B7A,
 16'hDD94, 16'h5061, 16'h2DA9, 16'hA94E,
 16'h97BA, 16'h5F3E, 16'h4FCA, 16'h9A2F,
 16'hDED7, 16'h5A24, 16'h33DF, 16'hB120,
 16'h86E0, 16'h4522, 16'h7FDA, 16'hE02A,
 16'h9AD1, 16'h1435, 16'h5EC5, 16'hDB42,
 16'hA2B7, 16'hE64E, 16'h54AD, 16'h5358,
 16'hA7A4, 16'h9A5F, 16'h539E, 16'h7B65,
 16'hC59A, 16'h8000, 16'h209B, 16'h6065,
 16'hD99C, 16'h9D63, 16'h049D, 16'h5A63,
 16'h239D, 16'hA464, 16'hCB9A, 16'h5968,
 16'h4395, 16'hA670, 16'hA48A, 16'h637D,
 16'h447A, 16'h9F90, 16'hD466, 16'h61A4,
 16'h1853, 16'h98B5, 16'h0243, 16'h50C5,
 16'h1734, 16'hA6D0, 16'hB02F, 16'h63D0,
 16'h2733, 16'hA7C6, 16'hC545, 16'h50AE,
 16'h7B62, 16'hA58A, 16'h968A, 16'h5562,
 16'h60B6, 16'hA22F, 16'h82ED, 16'h28F5,
 16'h722A, 16'hE6B8, 16'h9B64, 16'h1F82,
 16'h4D96, 16'h3054, 16'hAABF, 16'h8000,
 16'h50DA, 16'h781F, 16'hDBE2, 16'h9520,
 16'hF7DB, 16'h5E2F, 16'hF1C3, 16'h9F4F,
 16'h119A, 16'h5C81, 16'h0A61, 16'hB1C0,
 16'hB61D, 16'h4D07, 16'h7ED5, 16'hB650,
 16'h848B, 16'h3698, 16'h5646, 16'h03DB,
 16'hAE07, 16'h8515, 16'h54D0, 16'h7F48,
 16'hA9A3, 16'h9E6F, 16'h2B83, 16'h6788,
 16'h266F, 16'hA097, 16'hAC65, 16'h559D,
 16'h4964, 16'h9199, 16'hD56C, 16'h638D,
 16'hF07B, 16'hB17C, 16'hD48E, 16'h5569,
 16'h7B9F, 16'h9D59, 16'h9FAF, 16'h6548,
 16'h3CC3, 16'hA832, 16'h9FD8, 16'h3F1E,
 16'h7DEC, 16'hD30A, 16'h8D00, 16'h24F6,
 16'h5C13, 16'hC8E4, 16'hA325, 16'hEBD2,
 16'h5E37, 16'h4FC0, 16'hA249, 16'hBEAF,
 16'h5B59, 16'h549E, 16'hA36C, 16'h8D8B,
 16'h437E, 16'h6A7B, 16'h098A, 16'hAA72,
 16'h8092, 16'h486A, 16'h7F9B, 16'hAC61,
 16'hA2A1, 16'h1E5E, 16'h65A2, 16'h2060,
 16'h9E9D, 16'hD266, 16'h5C97, 16'h216C,
 16'hA991, 16'hB573, 16'h4D88, 16'h777E,
 16'hA67A, 16'h928E, 16'h316A, 16'h5F9E,
 16'h2A5B, 16'h9EAB, 16'h994D, 16'h61BC,
 16'h463C, 16'h9ECD, 16'hC72A, 16'h56DD,
 16'h6C1D, 16'hA5EA, 16'h8010, 16'h4DF7,
 16'h6D00, 16'hB409, 16'h9EEF, 16'h5818,
 16'h58E3, 16'hA220, 16'h95DF, 16'h5A22,
 16'h78DC, 16'hCA25, 16'h8FDC, 16'h1C24,
 16'h5DDD, 16'hBE20, 16'h9BE3, 16'h581A,
 16'h70EB, 16'hC410, 16'h90F5, 16'h0E05,
 16'h5C01, 16'hD8FA, 16'h930B, 16'h3EF0,
 16'h6315, 16'hD0E7, 16'hAA1C, 16'hD3E1,
 16'h4F21, 16'h7EDE, 16'hA324, 16'h8000,
 16'h3425, 16'h4EDC, 16'h1D22, 16'hA0E3,
 16'hB317, 16'h5EEE, 16'h340D, 16'hA5F7,
 16'hAA06, 16'h61FD, 16'h6601, 16'h9700,
 16'hBEFF, 16'h5E01, 16'h3C02, 16'hA7F9,
 16'h890D, 16'h4CEA, 16'h7F21, 16'hC1D3,
 16'hAD3B, 16'hEAB5, 16'h515C, 16'h7B92,
 16'h9A80, 16'h8002, 16'h55A7, 16'h6244,
 16'hD4D1, 16'h911A, 16'h0CFB, 16'h53F0,
 16'h0524, 16'hB1CA, 16'h9945, 16'h4EB0,
 16'h7FFF, 16'hBFA0, 16'hA865, 16'h5398,
 16'h5F68, 16'hA69B, 16'h9B60, 16'hF1A7,
 16'h5850, 16'h70BB, 16'h9C38, 16'h93D7,
 16'h6118, 16'h5FFA, 16'hB0F4, 16'h8A1F,
 16'h1BCE, 16'h6444, 16'hFBA9, 16'hAE6A,
 16'hF785, 16'h5B8B, 16'h2866, 16'h96A6,
 16'hF950, 16'h53BA, 16'h013D, 16'hADCB,
 16'h992E, 16'h4BD8, 16'h7F23, 16'hCCE0,
 16'h9D1F, 16'h29E1, 16'h4E1F, 16'hFBE0,
 16'hAE20, 16'h97E1, 16'h4A1F, 16'h7EDF,
 16'hBF23, 16'hA4DB, 16'h5026, 16'h5ADB,
 16'hAE23, 16'h90E0, 16'h261C, 16'h5EE9,
 16'hDB12, 16'hA2F2, 16'h330A, 16'h63FC,
 16'hC5FC, 16'hA90D, 16'h06EA, 16'h571F,
 16'h55D9, 16'h962E, 16'h93CB, 16'h663C,
 16'h3FBE, 16'h9C48, 16'hD2B2, 16'h5653,
 16'h3EA9, 16'h9E59, 16'h9FA7, 16'h6358,
 16'h4EAA, 16'h9E53, 16'hC6B0, 16'h654B,
 16'h28BC, 16'hA83D, 16'hBCCB, 16'h472C,
 16'h77DC, 16'hC61C, 16'h92ED, 16'h190A,
 16'h4D00, 16'hFAF6, 16'hAA13, 16'hCDE5,
 16'h5D22, 16'h40D9, 16'h962B, 16'hE7D3,
 16'h512D, 16'h28D5, 16'hAA27, 16'h85E0,
 16'h5716, 16'h75F5, 16'hB9FF, 16'hA90F,
 16'h4AE2, 16'h5A2E, 16'hADC0, 16'h9153,
 16'h3F99, 16'h5D7C, 16'hC86F, 16'hA9A5,
 16'h0648, 16'h63CA, 16'h1926, 16'hADE8,
 16'hCA0C, 16'h4AFE, 16'h70FA, 16'hBC0C,
 16'h8AF1, 16'h2E0F, 16'h47F6, 16'hAE01,
 16'hAB0A, 16'h15E9, 16'h6727, 16'h2BC7,
 16'hA74E, 16'hC89A, 16'h4F7F, 16'h6668,
 16'h9AB3, 16'h8A31, 16'h56EC, 16'h4AF6,
 16'hA627, 16'hACBF, 16'h595A, 16'h618E,
 16'h9E88, 16'h9E63, 16'h59AF, 16'h5142,
 16'hA4CB, 16'h992B, 16'h4ADB, 16'h5E21,
 16'h06E0, 16'hAC22, 16'hA2DA, 16'h622D,
 16'h55C9, 16'h9F43, 16'hC1B0, 16'h5C5E,
 16'h4294, 16'hA37A, 16'hAF77, 16'h459A,
 16'h6755, 16'hF2BB, 16'h9835, 16'hDCDB,
 16'h4517, 16'h29F6, 16'h9FFE, 16'hB60C,
 16'h63EB, 16'h331E, 16'hABDA, 16'hB82D,
 16'h45CD, 16'h6E37, 16'hFFC7, 16'hAC3A,
 16'hA6C6, 16'h5539, 16'h62C9, 16'h9735,
 16'hABCE, 16'h5A2F, 16'h53D4, 16'hAE28,
 16'h93DD, 16'h231E, 16'h5BE8, 16'hE812,
 16'hBCF3, 16'hE508, 16'h53FD, 16'h74FE,
 16'hAB07, 16'h99F4, 16'hEA10, 16'h48EC,
 16'h6C18, 16'h9DE3, 16'h8F22, 16'h54D9,
 16'h5A2C, 16'hB6D0, 16'hAE32, 16'hF9CD,
 16'h5634, 16'h4ACC, 16'h9833, 16'hC8CE,
 16'h5731, 16'h22D1, 16'hA52D, 16'hC1D5,
 16'h6028, 16'h2DDC, 16'hAA1F, 16'hC4E6,
 16'h4616, 16'h6AEF, 16'hDC0B, 16'hA9FA,
 16'hD402, 16'h4802, 16'h61FB, 16'h9B08,
 16'h96F4, 16'h540F, 16'h50F0, 16'hC110,
 16'hA5F1, 16'h170D, 16'h58F5, 16'hE208,
 16'hACFC, 16'h3BFF, 16'h5206, 16'hDDF6,
 16'hBD0D, 16'hC5F0, 16'h5213, 16'h71EA,
 16'hC119, 16'hAEE5, 16'hC91B, 16'h4AE7,
 16'h7715, 16'h9AF1, 16'hA609, 16'h10FD,
 16'h4DFB, 16'h5B0E, 16'h9DE9, 16'h9021,
 16'h1AD5, 16'h6033, 16'h17C5, 16'hAC43,
 16'hF3B6, 16'h4B51, 16'h30A8, 16'hA55C,
 16'h9BA2, 16'h465E, 16'h62A5, 16'hD256,
 16'hAEAF, 16'h194B, 16'h46BD, 16'hFB39,
 16'hABD3, 16'hE71F, 16'h5AEF, 16'h0203,
 16'hAA0B, 16'h28E7, 16'h4527, 16'hF7CB,
 16'hB443, 16'hA8B0, 16'h3C5A, 16'h6E9F,
 16'hD066, 16'hB098, 16'h3568, 16'h4D9A,
 16'hC462, 16'hACA4, 16'h2354, 16'h43B7,
 16'h263C, 16'hA2D3, 16'hA51B, 16'h62F9,
 16'h33F3, 16'hA921, 16'hDBCA, 16'h5D4B,
 16'h29A0, 16'hA974, 16'hE47A, 16'h5396,
 16'h2B5C, 16'hAEB0, 16'hA745, 16'h47C5,
 16'h5E33, 16'hB5D2, 16'hBB2C, 16'h0AD4,
 16'h592E, 16'h36CE, 16'h9A37, 16'hEAC2,
 16'h4848, 16'h02AC, 16'hB060, 16'hB193,
 16'h3B7A, 16'h6A7A, 16'hF293, 16'hAE5E,
 16'h08B1, 16'h4B41, 16'hD7CC, 16'hB128,
 16'h2DE2, 16'h4416, 16'hF6F2, 16'hB507,
 16'hC0FE, 16'h51FC, 16'h520A, 16'h9EF3,
 16'hA00E, 16'h41F2, 16'h560B, 16'hC7F9,
 16'hB303, 16'h4602, 16'h46F9, 16'hB20C,
 16'hAAEE, 16'h2718, 16'h4FE1, 16'hCF28,
 16'hB1CF, 16'h3C3B, 16'h4CBA, 16'hD550,
 16'hB0A6, 16'h0865, 16'h4092, 16'h2076,
 16'hAA81, 16'hA188, 16'h586F, 16'h5C9A,
 16'hCE5E, 16'hB7A8, 16'hE654, 16'h4EB0,
 16'h464C, 16'hA4B7, 16'hB046, 16'h5BBB,
 16'h3C47, 16'hA9B6, 16'hCB4E, 16'h55AD,
 16'h4558, 16'hA4A1, 16'hA568, 16'h378E,
 16'h577E, 16'hE375, 16'hBD98, 16'hD95A,
 16'h49B4, 16'h6A3F, 16'hAECE, 16'hA825,
 16'h26E8, 16'h460B, 16'hDE02, 16'hACF2,
 16'h3619, 16'h41DD, 16'hDA2C, 16'hBBCC,
 16'hC53B, 16'h55C0, 16'h5A43, 16'hABBB,
 16'hCD46, 16'h51BA, 16'h3C46, 16'hA0BB,
 16'hAD41, 16'h0AC4, 16'h5536, 16'h4CD2,
 16'hA426, 16'hB1E1, 16'h5917, 16'h3EF2,
 16'hAA06, 16'hAB02, 16'h38F5, 16'h5713,
 16'hD9E7, 16'hC51F, 16'hE3DC, 16'h4C28,
 16'h5BD4, 16'hA22E, 16'hBCD2, 16'h502D,
 16'h39D6, 16'hA925, 16'hA4E1, 16'h2818,
 16'h4DEF, 16'h000A, 16'hB8FD, 16'hF0FB,
 16'h4D0F, 16'h2BE6, 16'hA925, 16'hC3D1,
 16'h5C37, 16'h22C2, 16'hB245, 16'hD2B5,
 16'h4E51, 16'h56A9, 16'hB05C, 16'hA8A1,
 16'h225F, 16'h41A4, 16'hFC58, 16'hBDAC,
 16'hC64F, 16'h3DB6, 16'h6046, 16'hC0BF,
 16'hBB3B, 16'h4CC9, 16'h3834, 16'hA8CF,
 16'hB430, 16'h4FCF, 16'h4732, 16'hBCCC,
 16'hB138, 16'h10C3, 16'h4A43, 16'hEFB6,
 16'hBD52, 16'h12A5, 16'h4A65, 16'h0D90,
 16'hAF7C, 16'hE877, 16'h4C95, 16'h1260,
 16'hADA9, 16'hE350, 16'h4FB5, 16'h1B48,
 16'hAFB9, 16'hD847, 16'h4EB7, 16'h2F4D,
 16'hA1AE, 16'hE95A, 16'h4D9A, 16'hF375,
 16'hC07A, 16'hD498, 16'h4556, 16'h59BB,
 16'hBE34, 16'hBADE, 16'hFC10, 16'h4801,
 16'h32EE, 16'hA121, 16'hDBD2, 16'h4F39,
 16'h08BE, 16'hB149, 16'hEDB2, 16'h4251,
 16'h29AD, 16'hA853, 16'hBAAF, 16'h5B4E,
 16'h27B7, 16'hAF43, 16'hDCC4, 16'h4E33,
 16'h39D7, 16'hA720, 16'hB3E8, 16'h1512,
 16'h54F2, 16'h380B, 16'hA4F7, 16'hC208,
 16'h50F8, 16'h3F09, 16'hACF4, 16'hAA11,
 16'h49E8, 16'h3820, 16'hB1D7, 16'hC932,
 16'h04C6, 16'h6042, 16'h39B4, 16'hA357,
 16'hEFA0, 16'h3F68, 16'h1590, 16'hAD76,
 16'hA986, 16'h497E, 16'h4D80, 16'hC680,
 16'hBD80, 16'h207F, 16'h4184, 16'hF676,
 16'hBB93, 16'hE962, 16'h4EA9, 16'h2C4D,
 16'hADBC, 16'hC33B, 16'h4CCE, 16'h4329,
 16'hABE0, 16'hC817, 16'h4DF3, 16'h3503,
 16'hAC06, 16'hB0F1, 16'h3517, 16'h47E4,
 16'hEB20, 16'hC1DC, 16'hF427, 16'h45D6,
 16'h2E2E, 16'hAACE, 16'hB335, 16'h23CA,
 16'h5836, 16'hF8CA, 16'hB336, 16'h2EC9,
 16'h3339, 16'hD8C6, 16'hBD3A, 16'hDEC6,
 16'h523A, 16'h1DC6, 16'hB53A, 16'hE3C7,
 16'h4D37, 16'h39CC, 16'hA731, 16'hB2D1,
 16'h292D, 16'h4DD6, 16'hF727, 16'hC0DD,
 16'hD81E, 16'h36E6, 16'h5316, 16'hBAEE,
 16'hBC0F, 16'h47F3, 16'h300B, 16'hBAF7,
 16'hBD07, 16'hF3FB, 16'h4B04, 16'h3DFD,
 16'hA903, 16'hCAFC, 16'h5405, 16'h30FB,
 16'hAE06, 16'hBAF9, 16'h4508, 16'h43F6,
 16'hC10C, 16'hC3F3, 16'h240F, 16'h42EE,
 16'hE916, 16'hB8E5, 16'h2820, 16'h34DD,
 16'hD724, 16'hC1DB, 16'hED26, 16'h48D9,
 16'h3F29, 16'hA7D5, 16'hB32C, 16'h3FD2,
 16'h4230, 16'hF7D0, 16'hC02F, 16'hCFD2,
 16'h4D2D, 16'h4AD4, 16'hB22C, 16'hB5D3,
 16'h432D, 16'h35D2, 16'hCF30, 16'hC8CE,
 16'hE334, 16'h51C9, 16'h3E3A, 16'hB1C3,
 16'hD340, 16'h4ABC, 16'h4049, 16'hACB2,
 16'hB853, 16'h2DA8, 16'h3C5D, 16'hD59E,
 16'hC167, 16'h4393, 16'h3072, 16'hAD8C,
 16'hCF74, 16'h4F8D, 16'h2970, 16'hB094,
 16'hC468, 16'h409D, 16'h465C, 16'hE3AC,
 16'hC64B, 16'hD3C0, 16'h4A34, 16'h46D8,
 16'hAC1C, 16'hC0F1, 16'hFD02, 16'h4F0B,
 16'h34E8, 16'hB323, 16'hD0D4, 16'h4835,
 16'h3DC4, 16'hAF40, 16'hBBBD, 16'h2C44,
 16'h37BE, 16'hD440, 16'hC2C3, 16'h3C38,
 16'h38CF, 16'hD429, 16'hC0E0, 16'h1016,
 16'h42F5, 16'hEAFF, 16'hC90E, 16'hEEE5,
 16'h4228, 16'h4DCC, 16'hBC3F, 16'hBCB7,
 16'h1552, 16'h37A6, 16'hEF61, 16'hBB9A,
 16'h2769, 16'h3094, 16'hE86E, 16'hC492,
 16'hD06D, 16'h4D94, 16'h406A, 16'hB998,
 16'hCF67, 16'h469B, 16'h2D61, 16'hB6A5,
 16'hD354, 16'h0BB2, 16'h4D4A, 16'h2EB9,
 16'h9D45, 16'hAEBC, 16'h3543, 16'h37BE,
 16'hCE40, 16'hD2C3, 16'hE63A, 16'h42C8,
 16'h4C37, 16'hB5C9, 16'hC938, 16'hEAC7,
 16'h463A, 16'h3AC5, 16'hAF3C, 16'hCDC3,
 16'h103F, 16'h4CBE, 16'h0245, 16'hBBB9,
 16'hDE47, 16'h3CBA, 16'h4145, 16'hC1BB,
 16'hC145, 16'hF1BB, 16'h4444, 16'h17BE,
 16'hB43F, 16'h06C5, 16'h3638, 16'h08CA,
 16'hBA33, 16'hC3D1, 16'h4F2B, 16'h43DA,
 16'hCE20, 16'hC4E7, 16'h1A13, 16'h35F3,
 16'hDD07, 16'hC8FE, 16'h1CFE, 16'h3B07,
 16'hE7F4, 16'hCD11, 16'hE6EA, 16'h361A,
 16'h4EE3, 16'hC520, 16'hC7DE, 16'h4022,
 16'h29DF, 16'hC01E, 16'hBEE7, 16'h2615,
 16'h30EF, 16'hDA0C, 16'hD4FA, 16'hE8FF,
 16'h3C09, 16'h4BEE, 16'hC31B, 16'hCADD,
 16'h462B, 16'h2ACD, 16'hC039, 16'hCBC2,
 16'hE842, 16'h45BA, 16'h4B49, 16'hC0B5,
 16'hC94C, 16'hF8B6, 16'h3E45, 16'h30C1,
 16'hAB38, 16'hC7D0, 16'h1D28, 16'h44E1,
 16'h2715, 16'hB1F6, 16'hC0FD, 16'h4A11,
 16'h23E0, 16'hC22F, 16'hD7C4, 16'h1148,
 16'h51AD, 16'h0A5C, 16'hBE9D, 16'hDF69,
 16'h3792, 16'h3E72, 16'hC98B, 16'hC476,
 16'hEE8C, 16'h3F70, 16'h3795, 16'hAA63,
 16'hC6A7, 16'h494E, 16'h2BC0, 16'hB930,
 16'hD1E0, 16'h1510, 16'h4600, 16'h2DF0,
 16'hAF20, 16'hBFD0, 16'h3B40, 16'h33B1,
 16'hC75C, 16'hD698, 16'h4173, 16'h1E84,
 16'hB883, 16'hD178, 16'h438A, 16'h2C75,
 16'hBE8A, 16'hD179, 16'h3882, 16'h3285,
 16'hCB70, 16'hCA9D, 16'h1C54, 16'h37BC,
 16'hE834, 16'hC4DD, 16'h1411, 16'h3501,
 16'hE8EF, 16'hCA1F, 16'hF3D5, 16'h4036,
 16'h31BF, 16'hB24B, 16'hC7AE, 16'h2857,
 16'h36A7, 16'hE157, 16'hCBAD, 16'h0B4E,
 16'h31B9, 16'h163E, 16'hB2CC, 16'hDC29,
 16'h43E4, 16'h190E, 16'hB700, 16'hCFF1,
 16'h4320, 16'h36CE, 16'hC145, 16'hD6A8,
 16'h4369, 16'h1288, 16'hC285, 16'hD871,
 16'h2797, 16'h3E62, 16'hE8A3, 16'hCB59,
 16'hECAB, 16'h3E53, 16'h22AC, 16'hB457,
 16'hD2A4, 16'h3C63, 16'h3295, 16'hC274,
 16'hCF81, 16'hF48B, 16'h4268, 16'h3CA6,
 16'hB04C, 16'hC5C2, 16'h1630, 16'h38DD,
 16'hF417, 16'hC4F5, 16'h20FF, 16'h260D,
 16'hEAE8, 16'hCE22, 16'hD8D4, 16'h4434,
 16'h38C5, 16'hB942, 16'hD5B9, 16'h404A,
 16'h23B4, 16'hBE4C, 16'hD1B6, 16'h2948,
 16'h35BB, 16'hE041, 16'hCBC3, 16'h1D39,
 16'h29CC, 16'hF92F, 16'hC0D6, 16'hF224,
 16'h3CE3, 16'hF515, 16'hCDF3, 16'hEC07,
 16'h2AFE, 16'h44FD, 16'hF406, 16'hBBF8,
 16'hF30A, 16'h33F6, 16'hFD09, 16'hC6F8,
 16'hE105, 16'h3CFF, 16'h34FD, 16'hBC08,
 16'hD8F3, 16'h4312, 16'h21E9, 16'hBF1C,
 16'hCBDF, 16'h1526, 16'h37D5, 16'hF830,
 16'hC5CD, 16'h2234, 16'h27CC, 16'hD032,
 16'hD3D2, 16'h1B2A, 16'h37DA, 16'hE922,
 16'hCFE2, 16'hEE1A, 16'h2EEB, 16'h380F,
 16'hC3F9, 16'hD2FE, 16'h160B, 16'h30EC,
 16'h181B, 16'hB0E1, 16'hC722, 16'h3ADC,
 16'h2F25, 16'hDFDA, 16'hCF26, 16'hE0DC,
 16'h3821, 16'h34E2, 16'hC719, 16'hD3EF,
 16'h2A08, 16'h2B02, 16'hD5F3, 16'hD417,
 16'h02DF, 16'h402C, 16'h26C9, 16'hB442,
 16'hCCB4, 16'h2754, 16'h31A6, 16'hEF5F,
 16'hCA9D, 16'hDB67, 16'h3297, 16'h3968,
 16'hD69B, 16'hD160, 16'h0CA6, 16'h3354,
 16'hF1B4, 16'hD341, 16'hECCB, 16'h2D27,
 16'h3BE8, 16'hD50B, 16'hD200, 16'hEFF5,
 16'h3A15, 16'h29E3, 16'hB724, 16'hDAD7,
 16'h402B, 16'h22D6, 16'hBC26, 16'hCDDF,
 16'h1D1B, 16'h34EF, 16'hED05, 16'hD408,
 16'h09E9, 16'h3927, 16'h14C9, 16'hBD49,
 16'hD2A3, 16'h2B71, 16'h357C, 16'hF595,
 16'hC95C, 16'hD8B1, 16'h4042, 16'h2ECB,
 16'hC22B, 16'hD6DB, 16'hF723, 16'h3FDA,
 16'h332D, 16'hB4CB, 16'hD43F, 16'h28B4,
 16'h2D5C, 16'hDA92, 16'hD182, 16'h3468,
 16'h1BAE, 16'hD53C, 16'hD4DB, 16'hEF0E,
 16'h4108, 16'h23E2, 16'hC132, 16'hE2BC,
 16'h2D55, 16'h2F9C, 16'hEB70, 16'hC685,
 16'hE084, 16'h3A76, 16'h228E, 16'hC070,
 16'hE28E, 16'h3777, 16'h2382, 16'hC786,
 16'hDA70, 16'h389C, 16'h2557, 16'hC7B7,
 16'hD339, 16'h1BD7, 16'h2F19, 16'hFAF7,
 16'hC8FA, 16'hF414, 16'h3CDD, 16'h0532,
 16'hCFBF, 16'hF350, 16'h3BA2, 16'h1F6B,
 16'hBA89, 16'hD682, 16'h0475, 16'h4592,
 16'h1C68, 16'hBF9E, 16'hEC5D, 16'h36A7,
 16'h1C56, 16'hBAAC, 16'hD153, 16'h1DAD,
 16'h3155, 16'hF9A6, 16'hCA61, 16'hDC97,
 16'h1471, 16'h4288, 16'h0280, 16'hC477,
 16'hD694, 16'h1F5E, 16'h35B0, 16'hEA43,
 16'hCCCC, 16'hF925, 16'h32E9, 16'h0709,
 16'hCA04, 16'hEAF0, 16'h341C, 16'h1FD9,
 16'hC130, 16'hDAC8, 16'h293F, 16'h28BB,
 16'hE84B, 16'hCDAF, 16'hE356, 16'h32A7,
 16'h2D59, 16'hC8A9, 16'hDF55, 16'h38AD,
 16'h2050, 16'hC9B4, 16'hD947, 16'hFFBF,
 16'h363A, 16'h22CD, 16'hB92C, 16'hDCDC,
 16'h3E1C, 16'h1EEB, 16'hC60E, 16'hD5FA,
 16'h2EFE, 16'h1F09, 16'hD1F0, 16'hE217,
 16'h11E3, 16'h3A22, 16'h18DA, 16'hBF29,
 16'hD2D4, 16'h342E, 16'h25D1, 16'hD630,
 16'hD7D0, 16'h102E, 16'h2AD4, 16'hF92A,
 16'hD1DA, 16'hEA21, 16'h37E3, 16'h2418,
 16'hC9EF, 16'hDD0A, 16'h1CFE, 16'h2AF8,
 16'hE811, 16'hD3E8, 16'h0120, 16'h34D8,
 16'h142F, 16'hBFCA, 16'hDC3D, 16'h09BE,
 16'h4046, 16'h25B6, 16'hB74D, 16'hD6B1,
 16'h3850, 16'h17B0, 16'hC650, 16'hDCB1,
 16'h1F4C, 16'h2FB8, 16'hE942, 16'hD7C5,
 16'h1B34, 16'h1FD4, 16'hF223, 16'hCFE5,
 16'hFC13, 16'h34F7, 16'hF9FE, 16'hD20D,
 16'hFEE8, 16'h3323, 16'h15D4, 16'hC234,
 16'hD7C4, 16'h2D44, 16'h2AB5, 16'hD752,
 16'hDDA7, 16'h175F, 16'h2A9C, 16'h0569,
 16'hC492, 16'hEA73, 16'h3888, 16'h037D,
 16'hCC7F, 16'hE783, 16'h0C7C, 16'h4585,
 16'h087B, 16'hC984, 16'hFE7D, 16'h2782,
 16'h0380, 16'hC67D, 16'hD586, 16'h2378,
 16'h308A, 16'hE973, 16'hD892, 16'h0666,
 16'h2AA4, 16'h0551, 16'hC9BA, 16'hEA3D,
 16'h39CB, 16'h0F2C, 16'hCCDD, 16'hE91A,
 16'h2BF1, 16'h2604, 16'hCF05, 16'hD7F2,
 16'h0E18, 16'h29DF, 16'hFA2A, 16'hCFCD,
 16'hE939, 16'h11C3, 16'h3E41, 16'h06BC,
 16'hC747, 16'hDEB5, 16'h2E4E, 16'h1BB0,
 16'hC951, 16'hE1AF, 16'hFE51, 16'h39AE,
 16'h1F52, 16'hC0AF, 16'hDA50, 16'h0CB2,
 16'h324B, 16'h0AB5, 16'hCB4D, 16'hE4B1,
 16'h2D52, 16'h1BAB, 16'hCA57, 16'hE1A7,
 16'h1C5C, 16'h27A0, 16'hFB65, 16'hCA97,
 16'hF36D, 16'h2F8E, 16'h0F76, 16'hC486,
 16'hE580, 16'h387A, 16'h118B, 16'hCA71,
 16'hEA92, 16'h366B, 16'h1598, 16'hCA66,
 16'hE19A, 16'h1F68, 16'h2496, 16'hDF6B,
 16'hE094, 16'h266C, 16'h1A93, 16'hE470,
 16'hD28C, 16'h0B79, 16'h2681, 16'hE385,
 16'hE475, 16'hF691, 16'h1F69, 16'h329F,
 16'hDC57, 16'hDDB4, 16'h0241, 16'h2FCA,
 16'h1B2C, 16'hBEDD, 16'hD619, 16'h1CF2,
 16'h2403, 16'hE808, 16'hDBED, 16'h051D,
 16'h2EDA, 16'h0F2E, 16'hC7CA, 16'hE63E,
 16'h29BB, 16'h164B, 16'hD4B0, 16'hE353,
 16'h22AB, 16'h2556, 16'hE3AA, 16'hDB55,
 16'hEFAD, 16'h154F, 16'h38B6, 16'hF545,
 16'hCFC0, 16'h013B, 16'h21CA, 16'hEF30,
 16'hD6D7, 16'h0C22, 16'h23E4, 16'hEF17,
 16'hDBED, 16'h0E11, 16'h22F0, 16'h0010,
 16'hCDEE, 16'hF115, 16'h2FE7, 16'h0D1F,
 16'hCBDA, 16'hE22D, 16'h2CCB, 16'h223D,
 16'hE9BC, 16'hDB4C, 16'hF1AA, 16'h3360,
 16'h1396, 16'hCA75, 16'hE882, 16'h2384,
 16'h2277, 16'hE48D, 16'hD870, 16'h1192,
 16'h186E, 16'hE391, 16'hE370, 16'h088D,
 16'h3078, 16'hFF82, 16'hD586, 16'hF271,
 16'h0998, 16'h385E, 16'h08AD, 16'hC548,
 16'hDDC3, 16'h2333, 16'h1FD6, 16'hDD22,
 16'hE2E6, 16'hFA12, 16'h30F4, 16'h1C08,
 16'hC7FB, 16'hDE03, 16'h15FE, 16'h2401,
 16'hECFF, 16'hE002, 16'h07FC, 16'h2B06,
 16'h02F9, 16'hD209, 16'hE8F3, 16'h1311,
 16'h2EEA, 16'hE91C, 16'hDADF, 16'h1725,
 16'h15D7, 16'hE82C, 16'hDFD1, 16'hEB33,
 16'h11C8, 16'h383D, 16'hF5BF, 16'hD843,
 16'h0FBB, 16'h1847, 16'hEBB6, 16'hDF4F,
 16'hF6AC, 16'h3158, 16'h14A3, 16'hC862,
 16'hE59A, 16'hFC6B, 16'h2F8F, 16'h2577,
 16'hD384, 16'hE080, 16'h077E, 16'h2581,
 16'h0181, 16'hD07E, 16'hEB84, 16'h2B79,
 16'h168A, 16'hD271, 16'hE796, 16'h0D64,
 16'h29A2, 16'h0556, 16'hD2B4, 16'hE741,
 16'h15CA, 16'h2C2C, 16'h01DD, 16'hD11A,
 16'hE3F0, 16'h2905, 16'h1D07, 16'hE1EE,
 16'hE31A, 16'hF0DF, 16'h2927, 16'h1ED5,
 16'hD52E, 16'hEACF, 16'h1632, 16'h21CE,
 16'hF832, 16'hD6CF, 16'hF02F, 16'h2AD3,
 16'h172A, 16'hCCDA, 16'hE723, 16'h28E0,
 16'h101D, 16'hDCE5, 16'hE61A, 16'h0AE6,
 16'h321A, 16'hFBE6, 16'hDE1A, 16'hF2E6,
 16'h051A, 16'h34E4, 16'h061F, 16'hCCDE,
 16'hE625, 16'h21D7, 16'h192D, 16'hDCCF,
 16'hDF35, 16'hF1C9, 16'h2636, 16'h15CC,
 16'hD032, 16'hE8D0, 16'h112E, 16'h22D5,
 16'hF226, 16'hD9E1, 16'h1217, 16'h12F1,
 16'hE407, 16'hE502, 16'h02F4, 16'h2B16,
 16'h09DF, 16'hCF2C, 16'hEACA, 16'h0040,
 16'h31B7, 16'h1851, 16'hCDA8, 16'hDF5E,
 16'h069D, 16'h2366, 16'h0198, 16'hD66B,
 16'hF293, 16'h276E, 16'h0E92, 16'hD86A,
 16'hEB9C, 16'h1A5F, 16'h1DA5, 16'hF557,
 16'hD8AE, 16'hEC4B, 16'h29BE, 16'h1938,
 16'hD8D0, 16'hE62A, 16'h17DC, 16'h141F,
 16'hEFE5, 16'hE315, 16'hF0F2, 16'h2D0A,
 16'h11F9, 16'hDA04, 16'hECFD, 16'h0F02,
 16'h2A00, 16'hF900, 16'hD8FF, 16'hEC02,
 16'h0EFB, 16'h2B09, 16'h01F4, 16'hD20F,
 16'hEBED, 16'h2A16, 16'h0AE7, 16'hD01D,
 16'hEADE, 16'h0227, 16'h2CD5, 16'h1E2E,
 16'hD4CE, 16'hEA36, 16'hFEC7, 16'h293C,
 16'h18C2, 16'hD03E, 16'hE4C3, 16'h143C,
 16'h19C5, 16'hED3A, 16'hE3C7, 16'h0837,
 16'h1FCC, 16'hF932, 16'hDDD0, 16'hF52D,
 16'h22D5, 16'h132A, 16'hDCD8, 16'hE926,
 16'h10DB, 16'h2023, 16'hEDDF, 16'hE421,
 16'hF6DF, 16'h2021, 16'h1CDE, 16'hE022,
 16'hE6E0, 16'hF51F, 16'h27E1, 16'h131E,
 16'hD0E3, 16'hE91C, 16'h0AE7, 16'h2515,
 16'h07ED, 16'hD612, 16'hE6F0, 16'h1E0D,
 16'h19F7, 16'hE503, 16'hE904, 16'h12F5,
 16'h1C12, 16'hF2E6, 16'hE222, 16'hF3D6,
 16'h1C32, 16'h18C7, 16'hDB3F, 16'hEABB,
 16'h214B, 16'h10B0, 16'hDD55, 16'hECA7,
 16'hF45B, 16'h12A3, 16'h2E5F, 16'hE9A0,
 16'hEA61, 16'hF59E, 16'h0A61, 16'h27A2,
 16'hEB5A, 16'hDEAA, 16'h0951, 16'h14B5,
 16'hF446, 16'hDFBF, 16'hF23B, 16'h22CB,
 16'h142F, 16'hDCD9, 16'hEB1F, 16'h04E8,
 16'h2312, 16'h0AF3, 16'hD30A, 16'hE8F7,
 16'h200A, 16'h12F4, 16'hE00E, 16'hEDF0,
 16'h1912, 16'h11EB, 16'hE91A, 16'hE8E0,
 16'hF526, 16'h0CD3, 16'h2D36, 16'h04C0,
 16'hD44A, 16'hF0AC, 16'h235E, 16'h0398,
 16'hD672, 16'hEC84, 16'hFE85, 16'h2473,
 16'h1594, 16'hE065, 16'hECA2, 16'hFE58,
 16'h26AC, 16'h1151, 16'hD1B0, 16'hEB51,
 16'h12AE, 16'h0954, 16'hE7A8, 16'hEA5E,
 16'h199A, 16'h0F70, 16'hE884, 16'hEC8A,
 16'h0468, 16'h23A7, 16'h0249, 16'hE0C7,
 16'hF427, 16'h17ED, 16'h14FF, 16'hE614,
 16'hE9DA, 16'h0137, 16'h23B8, 16'h0958,
 16'hD299, 16'hE975, 16'h0C7F, 16'h208B,
 16'hFC6C, 16'hE09D, 16'hED5B, 16'h0CAC,
 16'h264F, 16'hF9B3, 16'hE44E, 16'hF4AF,
 16'h1A56, 16'h11A4, 16'hDD63, 16'hEC95,
 16'h0672, 16'h1F88, 16'h037E, 16'hD87B,
 16'hEB8E, 16'h0A68, 16'h24A2, 16'h0254,
 16'hDDB5, 16'hF644, 16'h1FC3, 16'h0936,
 16'hDAD1, 16'hEC28, 16'h09DE, 16'h1C1D,
 16'h01E7, 16'hE116, 16'hF1ED, 16'h200F,
 16'h0EF5, 16'hDB07, 16'hEFFD, 16'h15FF,
 16'h0D05, 16'hE5F6, 16'hED10, 16'h15EB,
 16'h1119, 16'hE7E2, 16'hEC23, 16'h15D8,
 16'h0E2E, 16'hECCC, 16'hEC38, 16'hFEC5,
 16'h233D, 16'h07C2, 16'hDB3F, 16'hEDC0,
 16'h0640, 16'h20C2, 16'h043C, 16'hDFC6,
 16'hF037, 16'h13CD, 16'h152E, 16'hEED8,
 16'hE521, 16'h01E7, 16'h1911, 16'hFCF7,
 16'hE300, 16'hF109, 16'h08F0, 16'h2815,
 16'h07E7, 16'hDA1D, 16'hEBDF, 16'h0F25,
 16'h17D7, 16'hF32B, 16'hE9D5, 16'hFD2A,
 16'h18D8, 16'h0A25, 16'hDCE0, 16'hFA1A,
 16'h19EC, 16'hFF0E, 16'hE2F8, 16'hFD03,
 16'h1E02, 16'hF6F8, 16'hE70F, 16'hF3EB,
 16'h0A1A, 16'h26E2, 16'hFA21, 16'hE0DD,
 16'hF326, 16'h14D8, 16'h1128, 16'hE8D9,
 16'hEC25, 16'h07DE, 16'h1220, 16'hF0E1,
 16'hED1D, 16'hF5E6, 16'h0516, 16'h2BEE,
 16'h050F, 16'hDCF3, 16'hED0B, 16'h0AF6,
 16'h160A, 16'hF0F5, 16'hEC0D, 16'h05F0,
 16'h1312, 16'hFFED, 16'hE114, 16'hEFEA,
 16'h171A, 16'h12E1, 16'hE924, 16'hF2D7,
 16'hFE2E, 16'h0DCF, 16'h1932, 16'hEACD,
 16'hEB33, 16'hF9CE, 16'h1430, 16'h12D3,
 16'hE529, 16'hEBDD, 16'h021B, 16'h18ED,
 16'hFF0B, 16'hE4FE, 16'hF7F9, 16'h1411,
 16'h0AE3, 16'hEA2B, 16'hF0C7, 16'hFF46,
 16'h1FAE, 16'h0B5D, 16'hE099, 16'hED70,
 16'h0788, 16'h187F, 16'hFA7C, 16'hE986,
 16'hFD79, 16'h1A87, 16'h097A, 16'hDE83,
 16'hEE81, 16'h0B7A, 16'h148D, 16'hFB6A,
 16'hE8A0, 16'hF754, 16'h17B9, 16'h0F3A,
 16'hE9D3, 16'hEE20, 16'h06ED, 16'h1205,
 16'hFA09, 16'hE8EA, 16'hF621, 16'h18D6,
 16'h0F32, 16'hEBC7, 16'hF13F, 16'hF3BC,
 16'h1148, 16'h10B7, 16'hE948, 16'hEEBA,
 16'hFC42, 16'h18C4, 16'h0736, 16'hDCD0,
 16'hF22A, 16'h15DC, 16'h061D, 16'hE5EB,
 16'hF50C, 16'hFBFE, 16'h13F9, 16'h160E,
 16'hECEB, 16'hF01B, 16'hFAE0, 16'h1725,
 16'h09D7, 16'hE02A, 16'hEFD7, 16'hFC27,
 16'h17DC, 16'h0E20, 16'hE8E5, 16'hF016,
 16'hFCF0, 16'h1A09, 16'h04FF, 16'hE5F8,
 16'hF413, 16'hFDE0, 16'h1A2E, 16'h10C5,
 16'hEC47, 16'hEEAE, 16'hF35C, 16'h0C9B,
 16'h166E, 16'hED89, 16'hF47F, 16'hF97A,
 16'h058C, 16'h1D6F, 16'hF396, 16'hEE66,
 16'h009E
};

logic [17:0] invader_depth;
logic invader_repeats;
assign invader_depth = 18'd3377; // same as numbers of samples
assign invader_repeats = 1;
/* end sine 441 hz*/

assign dout[15:0] = invader_ROM[adress][15:0];
assign repeats = invader_repeats;
assign depth = invader_depth;

endmodule 