// System-Verilog 'written by Alex Grinshpun May 2018
// New bitmap dudy February 2021
// (c) Technion IIT, Department of Electrical Engineering 2021 



module	alien_matrixBitMap	(	
					input	logic	clk,
					input	logic	resetN,
					input logic	[10:0] offsetX,// offset from top left  position 
					input logic	[10:0] offsetY,
					input	logic	InsideRectangle, //input that the pixel is within a bracket 
					input logic fireCollision, // if current alien was shot,
					input logic startOfFrame,
					input logic playGame, // wait for game to begin
					
					output	logic	drawingRequest, //output that the pixel should be dispalyed 
					output	logic	[7:0] RGBout,  //rgb value from the bitmap 
					output	logic	[3:0] HitEdgeCode, //one bit per edge 
					output	logic matrixDefeated,
					output	logic bottomAlien,
					output	logic [1:0] alienType



 ) ;

// this is the devider used to acess the right pixel 
localparam  int OBJECT_NUMBER_OF_Y_BITS = 5;  // 2^5 = 32 
localparam  int OBJECT_NUMBER_OF_X_BITS = 5;  // 2^5 = 32 

// never was read
/*const int ALIEN_WIDTH = 32;
const int ALIEN_HIGHT = 32;*/

localparam  int OBJECT_HEIGHT_Y = 1 <<  OBJECT_NUMBER_OF_Y_BITS ;
localparam  int OBJECT_WIDTH_X = 1 <<  OBJECT_NUMBER_OF_X_BITS;

// this is the devider used to acess the right pixel 
localparam  int OBJECT_HEIGHT_Y_DIVIDER = OBJECT_NUMBER_OF_Y_BITS - 2; //how many pixel bits are in every collision pixel
localparam  int OBJECT_WIDTH_X_DIVIDER =  OBJECT_NUMBER_OF_X_BITS - 2;

// generating a smiley bitmap


logic firstRow;
logic seconedRow;
logic thirdRow;
logic forthRow;

logic unsigned [0:3] [0:7] [0:1] initial_game   = 
	{{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
	{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1},
   {2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
	{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1}};

logic unsigned [0:3] [0:7] [0:1] MazeBiMapMask ;



logic [0:3] [0:OBJECT_HEIGHT_Y-1] [0:OBJECT_WIDTH_X-1] object_colors = {
{
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000011000000000110000000000,
	32'b00000000011000000000110000000000,
	32'b00000000011000000000110000000000,
	32'b00000000000110000011000000000000,
	32'b00000000000110000011000000000000,
	32'b00000000001110000011000000000000,
	32'b00000000011111111111110000000000,
	32'b00000000011111111111110000000000,
	32'b00000001111111111111111100000000,
	32'b00000001111001111100111100000000,
	32'b00000001111001111100111100000000,
	32'b00000011111111111111111110000000,
	32'b00000011111111111111111110000000,
	32'b00000011111111111111111110000000,
	32'b00000011111111111111111110000000,
	32'b00000011011111111111110110000000,
	32'b00000011011111111111110110000000,
	32'b00000011011000000000110110000000,
	32'b00000011011000000000110110000000,
	32'b00000011011111101111110110000000,
	32'b00000000000111101111000000000000,
	32'b00000000000111101111000000000000,
	32'b00000000000111101111000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000
	},
	
	
	{
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000001101100000000000000,
	32'b00000000000001101100000000000000,
	32'b00000000000001101100000000000000,
	32'b00000000000110000011000000000000,
	32'b00000000000110000011000000000000,
	32'b00000000001110000011000000000000,
	32'b00000000011111111111110000000000,
	32'b00000000011111111111110000000000,
	32'b00000001111111111111111100000000,
	32'b00000001111001111100111100000000,
	32'b00000001111001111100111100000000,
	32'b00000011111111111111111110000000,
	32'b00000011111111111111111110000000,
	32'b00000011111111111111111110000000,
	32'b00000011111111111111111110000000,
	32'b00000011011111111111110110000000,
	32'b00000011011111111111110110000000,
	32'b00000011011000000000110110000000,
	32'b00000011011000000000110110000000,
	32'b00000011011111101111110110000000,
	32'b00000000000110000011000000000000,
	32'b00000000000110000011000000000000,
	32'b00000000000110000011000000000000,
	32'b00000000011000000000110000000000,
	32'b00000000011000000000110000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000
	},
	
	{
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000111100000000000000,
	32'b00000000000000111100000000000000,
	32'b00000000000011111111000000000000,
	32'b00000000000011111111000000000000,
	32'b00000000000111111111100000000000,
	32'b00000000011111111111111000000000,
	32'b00000000011111111111111000000000,
	32'b00000001111100111100111110000000,
	32'b00000001111100111100111110000000,
	32'b00000001111111111111111110000000,
	32'b00000001111111111111111110000000,
	32'b00000000000011000011000000000000,
	32'b00000000000011000011000000000000,
	32'b00000000001100111100110000000000,
	32'b00000000011100111100111000000000,
	32'b00000000011100111100111000000000,
	32'b00000001100011000011001110000000,
	32'b00000001100011000011000110000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000
	},
	
	{
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000111100000000000000,
	32'b00000000000000111100000000000000,
	32'b00000000000011111111000000000000,
	32'b00000000000011111111000000000000,
	32'b00000000000111111111100000000000,
	32'b00000000011111111111111000000000,
	32'b00000000011111111111111000000000,
	32'b00000001111100111100111110000000,
	32'b00000001111100111100111110000000,
	32'b00000001111111111111111110000000,
	32'b00000001111111111111111110000000,
	32'b00000000001111111111110000000000,
	32'b00000000001100111100110000000000,
	32'b00000000001100111100110000000000,
	32'b00000000110000000000001100000000,
	32'b00000000110000000000001100000000,
	32'b00000000110000000000001100000000,
	32'b00000000001100000000110000000000,
	32'b00000000001100000000110000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000
	}

	};




//////////--------------------------------------------------------------------------------------------------------------=
//hit bit map has one bit per edge:  hit_colors[3:0] =   {Left, Top, Right, Bottom}	
//there is one bit per edge, in the corner two bits are set  



logic [0:3] [0:3] [3:0] hit_colors = 
		  {16'hC446,     
			16'h8C62,    
			16'h8932,
			16'h9113};

 

// pipeline (00) to get the pixel color from the array 	 

logic [6:0] frameCounter;

//////////--------------------------------------------------------------------------------------------------------------=
always_ff@(posedge clk or negedge playGame or negedge resetN)
begin
	if(!resetN || !playGame) begin
		MazeBiMapMask <= initial_game;
		frameCounter <= 0;
		matrixDefeated <= 0;

	end

	else begin
		
		if (startOfFrame) begin
			frameCounter <= frameCounter + 7'b1;
		end
	
		HitEdgeCode <= 4'h0;

		if ((InsideRectangle == 1'b1 )&(MazeBiMapMask[offsetY[8:5]][offsetX[8:5]] != 0 ))
		begin // inside an external bracket 
			HitEdgeCode <= hit_colors[offsetY >> OBJECT_HEIGHT_Y_DIVIDER][offsetX >> OBJECT_WIDTH_X_DIVIDER];	//get hitting edge from the colors table  
			if (fireCollision == 1) begin
				MazeBiMapMask[offsetY[8:5] ][offsetX[8:5]] <= 0; // to be replaced with explod
			end
			
		end 

		
		if (MazeBiMapMask == 0) begin
			MazeBiMapMask <= 
				{{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
				{2'd1,2'd1,2'd0,2'd1,2'd1,2'd1,2'd1,2'd1},
				{2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2,2'd2},
				{2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1,2'd1}};
			matrixDefeated <= 1;
		end
		else begin
			matrixDefeated <= 0;
		end
		
	end
		
end

//////////--------------------------------------------------------------------------------------------------------------=
// decide if to draw the pixel or not 
assign RGBout =	8'hFF;// white color
assign drawingRequest = (object_colors[frameCounter[6-2] + (2*((MazeBiMapMask[offsetY[8:5]][offsetX[8:5]]) -  1))][offsetY][offsetX] ) && InsideRectangle && playGame && MazeBiMapMask[offsetY[8:5] ][offsetX[8:5]]; // get optional transparent command from the bitmpap
always_comb begin
		if (offsetY[8:5] == 3'd3 && MazeBiMapMask[offsetY[8:5]][offsetX[8:5]] != 1'b0)begin
			 firstRow = 1'b1;
			 seconedRow = 1'b0;
			 thirdRow = 1'b0;
			 forthRow = 1'b0;
		end
		else if (offsetY[8:5] == 3'd2 && MazeBiMapMask[offsetY[8:5]][offsetX[8:5]] != 1'b0)begin
			 firstRow = 1'b0;
			 seconedRow = (MazeBiMapMask[3][offsetX[8:5]] == 1'b0) ? 1'b1 : 1'b0;
			 thirdRow = 1'b0;
			 forthRow = 1'b0;
			 
		end
		else if (offsetY[8:5] == 1'b1 && MazeBiMapMask[offsetY[8:5]][offsetX[8:5]] != 1'b0)begin
			 firstRow = 1'b0;
			 seconedRow = 1'b0;
			 thirdRow = ((MazeBiMapMask[3][offsetX[8:5]] == 1'b0) && (MazeBiMapMask[2][offsetX[8:5]] == 1'b0)) ? 1'b1 : 1'b0;
			 forthRow = 1'b0;
		end
		else if (offsetY[8:5] == 1'b0 && MazeBiMapMask[offsetY[8:5]][offsetX[8:5]] != 1'b0)begin
			firstRow = 1'b0;
			 seconedRow = 1'b0;
			 thirdRow = 1'b0;
			 forthRow = ((MazeBiMapMask[3][offsetX[8:5]] == 1'b0) && (MazeBiMapMask[2][offsetX[8:5]] == 1'b0) && (MazeBiMapMask[1][offsetX[8:5]] == 1'b0)) ? 1'b1 : 1'b0;
		end
		else begin
			 firstRow = 1'b0;
			 seconedRow = 1'b0;
			 thirdRow = 1'b0;
			 forthRow = 1'b0;		
			 end

		
end

assign bottomAlien =  (firstRow || seconedRow || thirdRow || forthRow) && drawingRequest;
assign alienType = MazeBiMapMask[offsetY[8:5]][offsetX[8:5]];

endmodule