module shot_ROM (
	
	input clk,
	input resetN,
	input [31:0] adress, // for future purpose
	output [15:0] dout,
	output [17:0] depth,
	output [31:0] repeats

);

/* shoot sound*/
 // stroe the value
bit [0:4079][15:0] shoot_ROM ={ // need to be 0 to 102 so first 2 bytes be on the left 
16'hFE3B, 16'hE468, 16'hE5E2, 16'h24F5,
 16'h5529, 16'h00BE, 16'h9E58, 16'hE894,
 16'h4B7D, 16'hF674, 16'hB69A, 16'hDB58,
 16'h0BB5, 16'h603E, 16'h17CE, 16'hBD27,
 16'hD2E3, 16'h1A14, 16'h37F5, 16'hE502,
 16'hCB06, 16'h00F3, 16'h5013, 16'h06EA,
 16'hAE18, 16'hDDE6, 16'hFC1C, 16'h4EE2,
 16'h251F, 16'hC7E2, 16'hCE1C, 16'h06E7,
 16'h4215, 16'hF4F0, 16'hC40A, 16'hF8FD,
 16'h4CFA, 16'h070F, 16'hBFE9, 16'hEA20,
 16'h0ED6, 16'h2C34, 16'hE8C1, 16'hB54A,
 16'hF9AB, 16'h4760, 16'h0496, 16'hCA73,
 16'hE885, 16'h5782, 16'h6A77, 16'hDB8F,
 16'hA96D, 16'hD495, 16'h226A, 16'hF296,
 16'hA16B, 16'hD094, 16'h156D, 16'h5090,
 16'h3774, 16'h4589, 16'h3E7A, 16'hF083,
 16'hDE7E, 16'h8C82, 16'h8000, 16'hCF83,
 16'h257B, 16'hEF89, 16'hF771, 16'h6E96,
 16'h7D63, 16'h7FA4, 16'hF455, 16'h80B2,
 16'h8000, 16'h80C0, 16'h8000, 16'h80C3,
 16'hD73F, 16'h6CBC, 16'h7D4C, 16'h7FAA,
 16'h7D65, 16'h7F86, 16'h3C92, 16'h8053,
 16'h8000, 16'h800D, 16'h931B, 16'h29B8,
 16'h2178, 16'h0757, 16'h7FDC, 16'h7CEF,
 16'h7FFF, 16'h3284, 16'hA6AF, 16'h8001,
 16'h8210, 16'h8CC2, 16'h826B, 16'hB96B,
 16'h28BB, 16'h7C23, 16'h7FFF, 16'h7BEA,
 16'h7FFF, 16'h7BBB, 16'hBE59, 16'h8000,
 16'h837A, 16'hA578, 16'hBE95, 16'hA85F,
 16'h03AD, 16'h4E48, 16'h7FFF, 16'h7A35,
 16'h7FFF, 16'h1228, 16'hB5DE, 16'h881D,
 16'h83E6, 16'h8000, 16'h8CE5, 16'h0420,
 16'h4CD7, 16'h4C35, 16'h6FBC, 16'h7A57,
 16'h7FFF, 16'h4C87, 16'h835B, 16'h8000,
 16'h8317, 16'h8B0E, 16'h92CD, 16'h9C59,
 16'h0180, 16'h7CA6, 16'h7FFC, 16'h7CEA,
 16'h7FFC, 16'h7A1A, 16'h11D5, 16'h8000,
 16'h81C2, 16'h8000, 16'hCDC0, 16'hC239,
 16'hCBD3, 16'h291D, 16'h7FFE, 16'h7CF3,
 16'h7FFE, 16'h66C5, 16'h0C51, 16'hB29B,
 16'h8276, 16'h8003, 16'h8A88, 16'hE777,
 16'hCF83, 16'hF88B, 16'h535F, 16'h7BBF,
 16'h7FFE, 16'h7C14, 16'h13B7, 16'hC185,
 16'h8837, 16'h8000, 16'h809E, 16'h8000,
 16'h06F5, 16'h2562, 16'h1E48, 16'h5B0D,
 16'h7D9E, 16'h7FB4, 16'h7CFD, 16'hD34F,
 16'h8000, 16'h82D7, 16'h8000, 16'h8345,
 16'h8000, 16'hD496, 16'h524C, 16'h63CB,
 16'h6125, 16'h7FFF, 16'h7B1A, 16'h7FFE,
 16'hEE28, 16'h83C8, 16'h8001, 16'h8393,
 16'hC78F, 16'hC149, 16'hABE5, 16'hFFE8,
 16'h4E50, 16'h7FFF, 16'h7CD0, 16'h7FE8,
 16'h5C63, 16'hF74E, 16'hB504, 16'h80AA,
 16'h8000, 16'h8007, 16'hF049, 16'h0369,
 16'hE7E1, 16'h36DA, 16'h7FFF, 16'h7D62,
 16'h7FFF, 16'h5B0D, 16'h0A0D, 16'hC6E5,
 16'h821D, 16'h8000, 16'h81F9, 16'hE42C,
 16'hE1A1, 16'hDFA0, 16'h3213, 16'h7D44,
 16'h7F5B, 16'h7E0F, 16'h7E81, 16'h3EF4,
 16'hF593, 16'h81E8, 16'h8001, 16'h82DE,
 16'hA8AB, 16'hFFC7, 16'hEFCE, 16'hFD93,
 16'h5917, 16'h7FFF, 16'h7990, 16'h7FFF,
 16'h6545, 16'hE7CA, 16'hAB35, 16'h85BD,
 16'h8000, 16'h8576, 16'h8AC3, 16'h05F8,
 16'h4A57, 16'h2852, 16'h3D0B, 16'h7FFF,
 16'h7AD5, 16'h7FFF, 16'h43AA, 16'h93EA,
 16'h8000, 16'h811B, 16'h8002, 16'h8062,
 16'hA7EE, 16'h19CA, 16'h4C75, 16'h3E57,
 16'h50D3, 16'h7E0C, 16'h7F0B, 16'h7DE9,
 16'h141A, 16'hC8EB, 16'h9407, 16'h8000,
 16'h80D5, 16'h8001, 16'hEF92, 16'h0B93,
 16'hF746, 16'h33E3, 16'h7EF5, 16'h7E30,
 16'h7EAE, 16'h6B70, 16'h5177, 16'hFA9E,
 16'h8000, 16'h80BA, 16'h8000, 16'hA1BA,
 16'hD350, 16'hD19F, 16'hF978, 16'h4F6C,
 16'h7DB4, 16'h7F28, 16'h7DFF, 16'h7ED8,
 16'h7F52, 16'h0283, 16'h80A7, 16'h8001,
 16'h80F7, 16'h9BE5, 16'h9F3A, 16'h9FAA,
 16'hF36D, 16'h3683, 16'h7F87, 16'h7D75,
 16'h7988, 16'h7D82, 16'h7F6D, 16'h60AA,
 16'hA239, 16'h8001, 16'h80ED, 16'h8000,
 16'hB78B, 16'hABAC, 16'hB91A, 16'h0022,
 16'h559F, 16'h7FA2, 16'h721D, 16'h7F23,
 16'h7D9F, 16'h7F9C, 16'h602A, 16'hA50F,
 16'h8003, 16'h8278, 16'h8000, 16'h8ECE,
 16'h9C10, 16'hE40D, 16'h26DB, 16'h6B38,
 16'h5CBB, 16'h674C, 16'h7AB3, 16'h7FFE,
 16'h7BC3, 16'h0F2E, 16'hA2E7, 16'h82FF,
 16'h8000, 16'h82BE, 16'h8000, 16'h8E6B,
 16'hDDC3, 16'h410C, 16'h3E27, 16'h2EA5,
 16'h7090, 16'h7FFF, 16'h7CFA, 16'h7FD3,
 16'h4D5E, 16'hB274, 16'h8004, 16'h8023,
 16'h8003, 16'h8000, 16'h8034, 16'hC5B7,
 16'h1459, 16'h679C, 16'h3F6A, 16'h3E96,
 16'h7766, 16'h7EA1, 16'h7F56, 16'h6AB3,
 16'h0C42, 16'hA6CC, 16'h8025, 16'h8000,
 16'h8005, 16'h8009, 16'h96EB, 16'hF61F,
 16'h4EDA, 16'h272B, 16'h22D2, 16'h5F2E,
 16'h7ED5, 16'h7E25, 16'h7EE4, 16'h5110,
 16'h07FE, 16'hBEF4, 16'h891A, 16'h8000,
 16'h8037, 16'h8000, 16'hD74C, 16'hF7AE,
 16'hF254, 16'h18AD, 16'h344F, 16'h7BB8,
 16'h7F3D, 16'h7DD2, 16'h641C, 16'h6DF9,
 16'h5AEF, 16'hD62C, 16'h8000, 16'h8068,
 16'h8000, 16'h80A6, 16'h943E, 16'hB6DE,
 16'h0106, 16'h4C14, 16'h46D3, 16'h3145,
 16'h6CA7, 16'h7F69, 16'h7D8A, 16'h677F,
 16'h4E7C, 16'h0987, 16'hC978, 16'h8187,
 16'h8002, 16'h8183, 16'h8002, 16'hDF7F,
 16'hE682, 16'hF17E, 16'h2F80, 16'h6283,
 16'h4979, 16'h588E, 16'h7D69, 16'h7FA1,
 16'h7D53, 16'h49BA, 16'hEE38, 16'hACD7,
 16'h8819, 16'h81F8, 16'h8000, 16'h8218,
 16'hD8DB, 16'hE62E, 16'hF0CE, 16'h2832,
 16'h53D2, 16'h7626, 16'h65E5, 16'h5A0B,
 16'h7D0B, 16'h7FDA, 16'h5F46, 16'h1696,
 16'hBD91, 16'h9745, 16'h8000, 16'h80E7,
 16'h8000, 16'hA783, 16'hE4B0, 16'hF01D,
 16'h0C14, 16'h44BD, 16'h5870, 16'h4467,
 16'h5BBC, 16'h7D25, 16'h7FF6, 16'h66F4,
 16'h351D, 16'h07D8, 16'hD12D, 16'h8FD3,
 16'h8127, 16'h8000, 16'h810D, 16'hBE06,
 16'hCEE2, 16'hEB39, 16'h19AB, 16'h4473,
 16'h706F, 16'h52AE, 16'h4F35, 16'h67E7,
 16'h7EFF, 16'h7E19, 16'h50D3, 16'h0F3C,
 16'hC6B8, 16'hA450, 16'h8000, 16'h8050,
 16'h8000, 16'h963F, 16'hE5D1, 16'hEA1C,
 16'h06FB, 16'h29EA, 16'h4833, 16'h77AE,
 16'h5D74, 16'h5368, 16'h69BC, 16'h7D20,
 16'h7FFF, 16'h41DE, 16'hF03E, 16'hA3A9,
 16'h866E, 16'h8001, 16'h8193, 16'h8000,
 16'h9BA6, 16'hFC59, 16'h00A3, 16'h0964,
 16'h2D90, 16'h3C81, 16'h606B, 16'h71AD,
 16'h5D37, 16'h54E7, 16'h69F9, 16'h7D29,
 16'h5DB5, 16'h0E6D, 16'hB671, 16'h81B0,
 16'h8030, 16'h8000, 16'h8001, 16'h8025,
 16'hC1C3, 16'h1A53, 16'h2F99, 16'h2178,
 16'h2B7A, 16'h2B92, 16'h5464, 16'h7AA4,
 16'h5C55, 16'h52B0, 16'h604E, 16'h73B3,
 16'h4A4C, 16'hFAB4, 16'hAE4D, 16'h89B2,
 16'h8150, 16'h80AD, 16'h8001, 16'h82A9,
 16'hCA58, 16'h19A8, 16'h2658, 16'h1FA8,
 16'h3058, 16'h4AA7, 16'h585A, 16'h43A6,
 16'h415A, 16'h5DA6, 16'h7759, 16'h6BA7,
 16'h3A5A, 16'h0FA3, 16'hE862, 16'hB499,
 16'h8000, 16'h808C, 16'h8001, 16'h8F7D,
 16'hBE8D, 16'hCE6B, 16'h049C, 16'h265C,
 16'h48AB, 16'h5750, 16'h2CB5, 16'h2047,
 16'h3DBC, 16'h7040, 16'h63C3, 16'h4D3C,
 16'h47C4, 16'h4E3F, 16'h4BBC, 16'hEC49,
 16'h93B1, 16'h8057, 16'h8000, 16'h8068,
 16'h8001, 16'h9280, 16'hD875, 16'h2397,
 16'h2D5D, 16'h22AC, 16'h274D, 16'h3ABA,
 16'h5740, 16'h36C4, 16'h2A3B, 16'h49C3,
 16'h5241, 16'h70B9, 16'h524F, 16'h2BA7,
 16'h1866, 16'hF189, 16'hC28C, 16'h805D,
 16'h8000, 16'h802B, 16'h8001, 16'h8EF2,
 16'hB52B, 16'hF2B8, 16'h1763, 16'h4784,
 16'h5595, 16'h3153, 16'h1DC3, 16'h2F29,
 16'h48E8, 16'h3F0B, 16'h3100, 16'h41F8,
 16'h5A0C, 16'h4EF3, 16'h290C, 16'h05F8,
 16'hD801, 16'hB509, 16'h82EA, 16'h8000,
 16'h80C9, 16'h8000, 16'hB6A0, 16'hCC77,
 16'hEB72, 16'h17A4, 16'h3446, 16'h52D0,
 16'h451B, 16'h25FA, 16'h28F1, 16'h3B23,
 16'h41CB, 16'h3545, 16'h38AE, 16'h4C5D,
 16'h599A, 16'h2D6E, 16'h148A, 16'h037D,
 16'hDA7E, 16'hBC85, 16'h8000, 16'h8086,
 16'h8000, 16'h8282, 16'hBF81, 16'hD77C,
 16'hEB87, 16'h1F76, 16'h448E, 16'h456D,
 16'h3398, 16'h2764, 16'h30A0, 16'h415B,
 16'h2CA9, 16'h1F53, 16'h36B2, 16'h3E49,
 16'h55BD, 16'h493A, 16'h1FD0, 16'h1827,
 16'h0BE0, 16'hE61A, 16'hA1EC, 16'h800D,
 16'h8000, 16'h81FB, 16'h860E, 16'h91E9,
 16'hC721, 16'hF2D5, 16'h2534, 16'h4BC4,
 16'h3744, 16'h29B4, 16'h3754, 16'h43A4,
 16'h2664, 16'h0F96, 16'h176D, 16'h3390,
 16'h4C74, 16'h4089, 16'h2E7A, 16'h3283,
 16'h397E, 16'h1C82, 16'h037E, 16'hDF83,
 16'hBB7C, 16'hA384, 16'h807C, 16'h8001,
 16'h807C, 16'h9684, 16'hCE7B, 16'hE784,
 16'hFD7E, 16'h1A80, 16'h3983, 16'h4979,
 16'h308B, 16'h2771, 16'h2793, 16'h3469,
 16'h299B, 16'h0D61, 16'h19A4, 16'h3357,
 16'h49AD, 16'h334F, 16'h27B4, 16'h274A,
 16'h2AB8, 16'h2946, 16'h00BB, 16'hD346,
 16'hACB7, 16'h9D4E, 16'h8FAB, 16'h8005,
 16'h829D, 16'h956B, 16'hBA8C, 16'hF67F,
 16'h0972, 16'h149F, 16'h2C50, 16'h2FC2,
 16'h422C, 16'h38E5, 16'h2409, 16'h1B09,
 16'h1BE6, 16'h292B, 16'h11C4, 16'h074C,
 16'h20A5, 16'h3869, 16'h3E8C, 16'h2B7D,
 16'h1B7C, 16'h2289, 16'h2774, 16'h0E8D,
 16'hEB76, 16'hD484, 16'hBB84, 16'h9072,
 16'h8003, 16'h875D, 16'h9CAE, 16'hB046,
 16'hB5C7, 16'hD52B, 16'hFFE4, 16'h2A0D,
 16'h3703, 16'h29ED, 16'h3222, 16'h39D1,
 16'h313A, 16'h1FBD, 16'h124A, 16'h16B1,
 16'h2053, 16'h10AB, 16'h0555, 16'h14AC,
 16'h2752, 16'h3BB1, 16'h294B, 16'h19BC,
 16'h1E3B, 16'h1ECE, 16'h1C28, 16'h01E3,
 16'hED13, 16'hDFF6, 16'hC401, 16'h9708,
 16'h84F1, 16'h8D15, 16'h96E5, 16'hB220,
 16'hC6DD, 16'hD024, 16'hE9DE, 16'h111E,
 16'h27E6, 16'h3B15, 16'h3EF2, 16'h2D06,
 16'h2A03, 16'h27F2, 16'h2D1A, 16'h20DB,
 16'h0A2E, 16'h0ACA, 16'h133D, 16'h0EBE,
 16'h0447, 16'h0CB4, 16'h1F4E, 16'h2FB2,
 16'h2D4D, 16'h1EB7, 16'h1942, 16'h14C6,
 16'h1330, 16'h15DD, 16'hFF15, 16'hECFA,
 16'hDAF4, 16'hB420, 16'hABCB, 16'hA14B,
 16'h8E9F, 16'h9776, 16'hA776, 16'hC59D,
 16'hD150, 16'hDFC2, 16'hFD2D, 16'h14E2,
 16'h3313, 16'h37F5, 16'h3105, 16'h2CFF,
 16'h2CFF, 16'h3101, 16'h2502, 16'h0FF8,
 16'h0F12, 16'h14E0, 16'h1530, 16'h09BF,
 16'hFD53, 16'h009B, 16'h0E77, 16'h1474,
 16'h18A3, 16'h1C47, 16'h21CE, 16'h281F,
 16'h13F1, 16'h0B00, 16'h070E, 16'h06E5,
 16'h0727, 16'hF5CF, 16'hE939, 16'hDBC1,
 16'hC942, 16'hADBE, 16'h9940, 16'h9EC5,
 16'hAC33, 16'hB5D7, 16'hBC1E, 16'hC9EE,
 16'hDB06, 16'hF606, 16'h11ED, 16'h1B21,
 16'h25D0, 16'h2D3F, 16'h35B3, 16'h375A,
 16'h279A, 16'h2170, 16'h1E87, 16'h1E81,
 16'h1B79, 16'h0D8B, 16'h0A72, 16'h0E8F,
 16'h0E72, 16'h038C, 16'hFF77, 16'h0184,
 16'h0A82, 16'h0F77, 16'h0892, 16'h0E64,
 16'h17A5, 16'h2252, 16'h1FB8, 16'h133E,
 16'h0ACD, 16'h0527, 16'h06E4, 16'h0113,
 16'hF2F5, 16'hF004, 16'hF502, 16'hEEFA,
 16'hD907, 16'hC2F9, 16'hB205, 16'hACFF,
 16'hB4FC, 16'hB40A, 16'hB9EF, 16'hC21A,
 16'hD3DB, 16'hE931, 16'hE7C2, 16'hF14C,
 16'h06A7, 16'h1C65, 16'h288F, 16'h2B7E,
 16'h2C75, 16'h2F98, 16'h305B, 16'h26B1,
 16'h1F45, 16'h18C3, 16'h1737, 16'h18CF,
 16'h0B2B, 16'h0ADA, 16'h0D23, 16'h0BDE,
 16'h0B23, 16'h01DA, 16'h032A, 16'h00D2,
 16'h0833, 16'h04C8, 16'hFF3D, 16'hFFBD,
 16'h0649, 16'h0BB1, 16'h0D55, 16'h0FA6,
 16'h115F, 16'h169B, 16'h106B, 16'h088F,
 16'h0175, 16'h008A, 16'hFD76, 16'h008A,
 16'hF277, 16'hEF86, 16'hF07F, 16'hF77B,
 16'hF68C, 16'hD66C, 16'hAD9C, 16'h8C5C,
 16'h8000, 16'h8646, 16'hB3C9, 16'hE025,
 16'h0AEF, 16'h1FFD, 16'h4817, 16'h7ED4,
 16'h7E42, 16'h2DA8, 16'hD16E, 16'hB97C,
 16'hB69A, 16'hE751, 16'h5BC2, 16'h4E2D,
 16'hD2E1, 16'hC614, 16'hC5F5, 16'hEF04,
 16'h6C00, 16'h49FF, 16'hD000, 16'hC404,
 16'hC7F4, 16'hF718, 16'h6ED8, 16'h4E3B,
 16'hCFB0, 16'hC267, 16'hC381, 16'hF498,
 16'h724D, 16'h4ACE, 16'hCE18, 16'hC002,
 16'hBFE6, 16'hF02F, 16'h70BE, 16'h4F52,
 16'hCDA1, 16'hBF69, 16'hBB91, 16'hEC72,
 16'h728E, 16'h526E, 16'hCC98, 16'hBA5E,
 16'hB7B1, 16'hE73D, 16'h73D7, 16'h5812,
 16'hD106, 16'hBAE1, 16'hBA39, 16'hE1AD,
 16'h686C, 16'h5F7B, 16'hD29D, 16'hB34E,
 16'hBAC4, 16'hD62D, 16'h5DDF, 16'h6B18,
 16'hE1ED, 16'hB413, 16'hB9E8, 16'hD022,
 16'h4CD0, 16'h7941, 16'hF5AB, 16'hB26D,
 16'hB676, 16'hC7AB, 16'h3632, 16'h7EF3,
 16'h09E7, 16'hB33E, 16'hB89E, 16'hBE86,
 16'h2657, 16'h7ECA, 16'h2317, 16'hB706,
 16'hB4E1, 16'hB932, 16'h0DC1, 16'h7F45,
 16'h3DBC, 16'hBB3D, 16'hB2D0, 16'hB81D,
 16'hF1FA, 16'h7FEB, 16'h5435, 16'hCBA6,
 16'hB285, 16'hB64B, 16'hDFE9, 16'h66E1,
 16'h7355, 16'hDF75, 16'hABC2, 16'hB508,
 16'hCE2B, 16'h46A5, 16'h7FFF, 16'h0353,
 16'hAFCE, 16'hB717, 16'hBFFE, 16'h20F4,
 16'h7FFF, 16'h2EF0, 16'hB608, 16'hB508,
 16'hB8E1, 16'hF73D, 16'h7FFF, 16'h548F,
 16'hC140, 16'hADF5, 16'hB2D4, 16'hE165,
 16'h6D5F, 16'h74DE, 16'hE0E6, 16'hAE55,
 16'hBA72, 16'hCBC3, 16'h3D0D, 16'h7FFF,
 16'h13BD, 16'hAF62, 16'hB284, 16'hB891,
 16'h0C60, 16'h7FA9, 16'h4753, 16'hBAAB,
 16'hAE5C, 16'hB298, 16'hE378, 16'h7374,
 16'h71A4, 16'hDB41, 16'hAADC, 16'hB305,
 16'hC51A, 16'h3DC8, 16'h7E55, 16'h1791,
 16'hAD87, 16'hB562, 16'hB9B3, 16'h003A,
 16'h7ED8, 16'h531A, 16'hC3F0, 16'hAB09,
 16'hB1FB, 16'hDB03, 16'h5DFE, 16'h7F02,
 16'hF3FE, 16'hAA03, 16'hB5FA, 16'hBC0A,
 16'h23F1, 16'h7E13, 16'h3AEC, 16'hB313,
 16'hACEF, 16'hB50E, 16'hE5F4, 16'h780B,
 16'h75F8, 16'hDD03, 16'hA902, 16'hB5F8,
 16'hC010, 16'h2FE9, 16'h7E1E, 16'h2DDA,
 16'hAF2D, 16'hACCD, 16'hB63A, 16'hEFC0,
 16'h7F44, 16'h6AB8, 16'hD14A, 16'hA6B7,
 16'hB648, 16'hC6B9, 16'h3144, 16'h7EC0,
 16'h273B, 16'hAECB, 16'hAF2F, 16'hB9D7,
 16'hEE24, 16'h7BE1, 16'h7518, 16'hD7EF,
 16'hAE0A, 16'hB1FF, 16'hC6F8, 16'h3010,
 16'h7DE7, 16'h3422, 16'hB1D7, 16'hAD2F,
 16'hB5CA, 16'hE43D, 16'h6ABC, 16'h7E4B,
 16'hE9AF, 16'hA856, 16'hB5A5, 16'hC060,
 16'h179C, 16'h7E68, 16'h4E94, 16'hBE6F,
 16'hA68F, 16'hB273, 16'hD78C, 16'h4975,
 16'h7E89, 16'h0B79, 16'hA786, 16'hAF7B,
 16'hB685, 16'hF77A, 16'h7E87, 16'h7079,
 16'hD087, 16'hA87B, 16'hB381, 16'hC484,
 16'h2177, 16'h7F8E, 16'h3D6D, 16'hB398,
 16'hAC63, 16'hB2A3, 16'hDC57, 16'h56AD,
 16'h7E50, 16'h07B4, 16'hA748, 16'hB4BC,
 16'hB83F, 16'hF7C4, 16'h7E3D, 16'h71C0,
 16'hD745, 16'hA8B3, 16'hB555, 16'hC5A3,
 16'h1B67, 16'h7F8D, 16'h4E81, 16'hBB6E,
 16'hAAA5, 16'hB447, 16'hD4CF, 16'h3D1A,
 16'h7EFD, 16'h24EC, 16'hAE2A, 16'hAEC2,
 16'hBB51, 16'hE49D, 16'h5D72, 16'h7E82,
 16'hFC89, 16'hA86D, 16'hB09A, 16'hBB63,
 16'hFA9D, 16'h7D67, 16'h7391, 16'hDE79,
 16'hA57C, 16'hB192, 16'hC65E, 16'h0FB3,
 16'h7E39, 16'h5CDC, 16'hC210, 16'hA905,
 16'hB5E6, 16'hCA2C, 16'h23C4, 16'h7E4B,
 16'h47A8, 16'hB663, 16'hAA95, 16'hB46F,
 16'hD391, 16'h376C, 16'h7E9A, 16'h305E,
 16'hB1AD, 16'hAD44, 16'hB8CE, 16'hDE1E,
 16'h48F8, 16'h7DF2, 16'h1C24, 16'hAEC4,
 16'hAE55, 16'hBB92, 16'hE486, 16'h5764,
 16'h7FAE, 16'h0944, 16'hACC8, 16'hB02F,
 16'hBDD6, 16'hEF27, 16'h5FDA, 16'h7E2A,
 16'hFDCE, 16'hAB3D, 16'hB2B3, 16'hC060,
 16'hF08C, 16'h648A, 16'h7E5E, 16'hF8BB,
 16'hA72A, 16'hAEF1, 16'hBEF6, 16'hF322,
 16'h6AC7, 16'h7F4E, 16'hF79F, 16'hAE72,
 16'hAF81, 16'hBF88, 16'hF671, 16'h6693,
 16'h7E6D, 16'hF590, 16'hAA77, 16'hB17E,
 16'hC390, 16'hF35F, 16'h64B6, 16'h7E32,
 16'hFFE7, 16'hAE01, 16'hAE17, 16'hC2D1,
 16'hEF47, 16'h5AA0, 16'h7E79, 16'h0671,
 16'hAFA2, 16'hB34E, 16'hBFBF, 16'hEB38,
 16'h4CCF, 16'h7E2C, 16'h19D5, 16'hB12D,
 16'hAFCF, 16'hBC39, 16'hE1BB, 16'h3F52,
 16'h7E9E, 16'h2975, 16'hB178, 16'hB19A,
 16'hBA53, 16'hDAC0, 16'h2D2D, 16'h7DE6,
 16'h4308, 16'hB907, 16'hA5EE, 16'hAE1B,
 16'hCBDC, 16'h152C, 16'h7DCE, 16'h5036,
 16'hBFCA, 16'hA232, 16'hB1D4, 16'hCE24,
 16'h07E6, 16'h7F0F, 16'h68FC, 16'hCEF8,
 16'hA815, 16'hB1DE, 16'hC730, 16'hF6C2,
 16'h684B, 16'h7DA9, 16'hF062, 16'hAA94,
 16'hAE75, 16'hC283, 16'hE984, 16'h4876,
 16'h7F8E, 16'h1E6F, 16'hAF94, 16'hAD6A,
 16'hBC96, 16'hDA6B, 16'h2A94, 16'h7E6E,
 16'h4790, 16'hBE71, 16'hAD8E, 16'hB672,
 16'hD28F, 16'h0C70, 16'h7F90, 16'h7170,
 16'hDA90, 16'hAF6F, 16'hB193, 16'hCA6B,
 16'hF597, 16'h5367, 16'h7F9A, 16'h1166,
 16'hAF9A, 16'hAE66, 16'hBE9A, 16'hE467,
 16'h2697, 16'h7E6D, 16'h498C, 16'hBE7D,
 16'hAF79, 16'hB792, 16'hD462, 16'h06AB,
 16'h7347, 16'h7CC8, 16'hE927, 16'hABEA,
 16'hB705, 16'hC60C, 16'hEEE4, 16'h3C2A,
 16'h7DC9, 16'h3142, 16'hB5B6, 16'hAF4F,
 16'hB6AF, 16'hDA50, 16'h11B4, 16'h7B44,
 16'h72C8, 16'hDB26, 16'hAEF2, 16'hB5F1,
 16'hCC30, 16'hF0AD, 16'h3E77, 16'h7E63,
 16'h27C4, 16'hB516, 16'hB010, 16'hBDCA,
 16'hDD5B, 16'h0E81, 16'h7AA1, 16'h7141,
 16'hE0D7, 16'hB118, 16'hB3F2, 16'hC80B,
 16'hEAF1, 16'h361A, 16'h7FD3, 16'h3748,
 16'hB995, 16'hAE96, 16'hB638, 16'hD5FE,
 16'h05C8, 16'h6776, 16'h7F48, 16'hF2FE,
 16'hB1BA, 16'hB38E, 16'hBF2D, 16'hEA13,
 16'h21B2, 16'h7FFD, 16'h5448, 16'hC3E3,
 16'hADFA, 16'hB620, 16'hD1D0, 16'hF836,
 16'h45CD, 16'h7FFF, 16'h1DF3, 16'hB7EB,
 16'hB13F, 16'hBB8E, 16'hDDAD, 16'h0C13,
 16'h7133, 16'h7B81, 16'hEBCE, 16'hAFE2,
 16'hB26F, 16'hC241, 16'hE50C, 16'h1DA9,
 16'h7F9E, 16'h5620, 16'hC81D, 16'hAFAD,
 16'hB381, 16'hCE58, 16'hF3C7, 16'h3022,
 16'h7FFF, 16'h3709, 16'hBBF7, 16'hAC12,
 16'hB6DE, 16'hD539, 16'hFCAA, 16'h4976,
 16'h7FFF, 16'h16C3, 16'hB310, 16'hAE20,
 16'hBDAD, 16'hDE87, 16'h0746, 16'h60ED,
 16'h7EDF, 16'hFA55, 16'hB277, 16'hB4BD,
 16'hC012, 16'hE21B, 16'h0EB9, 16'h7272,
 16'h6E66, 16'hE6C0, 16'hAE1C, 16'hB104,
 16'hC5DF, 16'hE83D, 16'h10A9, 16'h7F6F,
 16'h667B, 16'hD499, 16'hB054, 16'hB5BD,
 16'hC835, 16'hE7D7, 16'h1A20, 16'h7FE6,
 16'h5C16, 16'hD4EC, 16'hB114, 16'hB6EC,
 16'hCD16, 16'hEAE6, 16'h1D1F, 16'h7FDA,
 16'h5E30, 16'hCEC5, 16'hB347, 16'hB7AB,
 16'hC864, 16'hEB8D, 16'h1882, 16'h7F6E,
 16'h60A3, 16'hD54C, 16'hB1C4, 16'hB72D,
 16'hC9E1, 16'hEA12, 16'h15FA, 16'h7FFB,
 16'h630F, 16'hD8E9, 16'hB21E, 16'hB5DB,
 16'hC92B, 16'hE9D0, 16'h1235, 16'h74C6,
 16'h6D3E, 16'hE9BE, 16'hB147, 16'hB1B3,
 16'hC954, 16'hE6A2, 16'h0A6A, 16'h6689,
 16'h7986, 16'hFD69, 16'hB4A9, 16'hB543,
 16'hBFD4, 16'hE513, 16'h0008, 16'h4FDB,
 16'h7E43, 16'h129D, 16'hB685, 16'hB359,
 16'hBDC8, 16'hD918, 16'hF907, 16'h3DDB,
 16'h7FFC, 16'h2EA2, 16'hBE78, 16'hAC72,
 16'hBA9F, 16'hD556, 16'hF3B0, 16'h224E,
 16'h7FAE, 16'h515B, 16'hC797, 16'hB47D,
 16'hB56A, 16'hCCB3, 16'hEE2B, 16'h10FB,
 16'h72DB, 16'h6F53, 16'hEB7E, 16'hB6B1,
 16'hB61F, 16'hC111, 16'hE7BF, 16'h0071,
 16'h4861, 16'h7FCA, 16'h1B0E, 16'hBA16,
 16'hB1CC, 16'hBA4C, 16'hE0A1, 16'hF46D,
 16'h288B, 16'h7FFF, 16'h4D8E, 16'hCB67,
 16'hB0AA, 16'hB63F, 16'hCCDC, 16'hF105,
 16'h0D1F, 16'h64BA, 16'h7B6F, 16'h0067,
 16'hB5C3, 16'hB313, 16'hBF16, 16'hE5C3,
 16'hFA63, 16'h3379, 16'h7FA6, 16'h413F,
 16'hC3DA, 16'hAE11, 16'hB9FE, 16'hD6F7,
 16'hF010, 16'h0DF0, 16'h690B, 16'h77FC,
 16'hFAF9, 16'hB915, 16'hB7DB, 16'hC237,
 16'hE6B4, 16'hF564, 16'h3082, 16'h7D98,
 16'h434F, 16'hC6C9, 16'hB321, 16'hB9F4,
 16'hD2F7, 16'hF01C, 16'h06D4, 16'h583B,
 16'h7DB8, 16'h1652, 16'hB5A6, 16'hB35F,
 16'hBB9F, 16'hDB62, 16'hF29E, 16'h1E61,
 16'h7CA1, 16'h645B, 16'hE2AB, 16'hB54D,
 16'hB9BC, 16'hC73A, 16'hE6D1, 16'hFA24,
 16'h31E6, 16'h7F11, 16'h41F7, 16'hC402,
 16'hB405, 16'hBBF4, 16'hD013, 16'hF0E6,
 16'h0720, 16'h4EDB, 16'h7E2A, 16'h23D2,
 16'hBD31, 16'hB1CB, 16'hBA38, 16'hD7C7,
 16'hF73A, 16'h0EC6, 16'h6138, 16'h7DC9,
 16'h0936, 16'hB8CD, 16'hB630, 16'hBED3,
 16'hDE29, 16'hF6DC, 16'h191F, 16'h6EE6,
 16'h6F16, 16'hEFEE, 16'hB50E, 16'hB9F6,
 16'hC406, 16'hE700, 16'hF6FA, 16'h1B0B,
 16'h75F0, 16'h5F15, 16'hDFE7, 16'hAE1D,
 16'hAEDE, 16'hC128, 16'hE3D2, 16'hF633,
 16'h1DC8, 16'h753D, 16'h5FBE, 16'hDD48,
 16'hB1B1, 16'hB755, 16'hC0A7, 16'hE95D,
 16'hF99E, 16'h1E66, 16'h7795, 16'h5C71,
 16'hE28A, 16'hB37B, 16'hB67F, 16'hC385,
 16'hE879, 16'hFD88, 16'h1B78, 16'h7388,
 16'h6377, 16'hEC8B, 16'hB673, 16'hB28F,
 16'hC56F, 16'hE492, 16'hF96E, 16'h1992,
 16'h666E, 16'h7192, 16'hFF6E, 16'hB692,
 16'hB66E, 16'hC092, 16'hE16D, 16'hF794,
 16'h0F6C, 16'h5794, 16'h7E6B, 16'h1896,
 16'hBA68, 16'hB69A, 16'hBD65, 16'hDB9D,
 16'hF560, 16'h08A3, 16'h415B, 16'h7FA6,
 16'h345A, 16'hC0A6, 16'hB259, 16'hBEA9,
 16'hD455, 16'hECAD, 16'hFD52, 16'h2BAE,
 16'h7E52, 16'h59AE, 16'hDD53, 16'hB8AC,
 16'hB955, 16'hC6A9, 16'hEB5A, 16'hF9A3,
 16'h1760, 16'h619C, 16'h7369, 16'h0C92,
 16'hB774, 16'hB385, 16'hC281, 16'hDD7A,
 16'hF58B, 16'h0770, 16'h3A95, 16'h7F66,
 16'h3E9F, 16'hCA5C, 16'hB3A8, 16'hBA54,
 16'hD1B0, 16'hEC4D, 16'hFDB6, 16'h1947,
 16'h64BB, 16'h7543, 16'h01C0, 16'hB83D,
 16'hB8C5, 16'hC33A, 16'hDEC7, 16'hF639,
 16'h03C6, 16'h363A, 16'h7EC7, 16'h4438,
 16'hCCC9, 16'hB537, 16'hBBC8, 16'hCE39,
 16'hE8C6, 16'hFD3B, 16'h14C4, 16'h563D,
 16'h7DC1, 16'h1942, 16'hBBBC, 16'hB545,
 16'hBEB9, 16'hD749, 16'hF3B5, 16'hFE4E,
 16'h24AF, 16'h7253, 16'h60AB, 16'hF056,
 16'hB8A9, 16'hB25A, 16'hC1A3, 16'hE05F,
 16'hF69E, 16'h0864, 16'h339C, 16'h7F64,
 16'h499D, 16'hCE60, 16'hB5A3, 16'hB659,
 16'hC6AC, 16'hE54F, 16'hF9B7, 16'h0D41,
 16'h42C7, 16'h7E31, 16'h34D9, 16'hC31D,
 16'hB4EC, 16'hBB0A, 16'hCE00, 16'hEBF7,
 16'hFC13, 16'h0FE2, 16'h4629, 16'h7DCD,
 16'h2B3B, 16'hC1BF, 16'hB247, 16'hB7B3,
 16'hD454, 16'hEBA5, 16'hFD5F, 16'h0FA0,
 16'h4960, 16'h7EA1, 16'h285E, 16'hC0A3,
 16'hB15B, 16'hB9A8, 16'hD453, 16'hEFB4,
 16'hFF46, 16'h11C0, 16'h4539, 16'h7BCE,
 16'h2D2A, 16'hC2E0, 16'hB216, 16'hB8F4,
 16'hD103, 16'hE904, 16'hFAF6, 16'h0A10,
 16'h3DEB, 16'h7C1A, 16'h38E0, 16'hC725,
 16'hB1D7, 16'hB92D, 16'hCECF, 16'hEC34,
 16'hFCCA, 16'h0937, 16'h2FC9, 16'h7836,
 16'h4ECB, 16'hDB35, 16'hB9CB, 16'hBB34,
 16'hC7CD, 16'hE332, 16'hF5D0, 16'h052E,
 16'h1FD4, 16'h6528, 16'h6ADD, 16'h011E,
 16'hB9E7, 16'hB314, 16'hC1F0, 16'hDE0C,
 16'hEFF9, 16'hFE02, 16'h1203, 16'h45F7,
 16'h7B0F, 16'h2DEB, 16'hC21B, 16'hB1E0,
 16'hBC26, 16'hD3D4, 16'hE931, 16'hFFC9,
 16'h083E, 16'h23BC, 16'h734A, 16'h5AB0,
 16'hE756, 16'hB8A3, 16'hB564, 16'hC195,
 16'hE071, 16'hF28B, 16'h0278, 16'h1086,
 16'h467B, 16'h7785, 16'h2A7A, 16'hC287,
 16'hB179, 16'hBC88, 16'hCE76, 16'hEE8C,
 16'hFD71, 16'h0493, 16'h2268, 16'h669E,
 16'h645B, 16'hFCAD, 16'hBA4B, 16'hB0BC,
 16'hC03C, 16'hDDCE, 16'hF028, 16'hFFE2,
 16'h0C13, 16'h30F6, 16'h7802, 16'h4A07,
 16'hDBF0, 16'hBA19, 16'hB4DE, 16'hC82A,
 16'hE2CF, 16'hF537, 16'h03C4, 16'h1241,
 16'h3DBB, 16'h7846, 16'h3ABB, 16'hCA44,
 16'hB4BE, 16'hB83E, 16'hD0C6, 16'hE935,
 16'hF5D2, 16'h0427, 16'h0FE0, 16'h4718,
 16'h7EF1, 16'h3005, 16'hC206, 16'hB5EF,
 16'hBC1B, 16'hCFDC, 16'hED2C, 16'hFACE,
 16'h0838, 16'h0EC1, 16'h4445, 16'h7BB7,
 16'h2C4D, 16'hC6B0, 16'hB551, 16'hBAAF,
 16'hD151, 16'hE9B1, 16'hF64B, 16'h08BA,
 16'h0F40, 16'h3DC7, 16'h7A33, 16'h3AD3,
 16'hCD26, 16'hB4E1, 16'hBF18, 16'hCBF0,
 16'hE608, 16'hF5FE, 16'h04FC, 16'h0F0A,
 16'h30F2, 16'h6F10, 16'h49EF, 16'hE210,
 16'hB5F3, 16'hB50A, 16'hC9FA, 16'hE201,
 16'hF604, 16'h02F8, 16'h090C, 16'h22EF,
 16'h6018, 16'h66DF, 16'h042A, 16'hBBCE,
 16'hB038, 16'hBEC4, 16'hDE3F, 16'hF1BF,
 16'hFE42, 16'h0BBE, 16'h1840, 16'h42C3,
 16'h783A, 16'h31CB, 16'hC72E, 16'hB6DA,
 16'hB61B, 16'hCDF2, 16'hEC01, 16'hF70C,
 16'h05E7, 16'h1026, 16'h26CD, 16'h6140,
 16'h62B3, 16'h015A, 16'hBD9A, 16'hB271,
 16'hBD86, 16'hDB82, 16'hEF78, 16'h008C,
 16'h0A71, 16'h1090, 16'h3B71, 16'h6F8D,
 16'h4676, 16'hDC85, 16'hBA81, 16'hB978,
 16'hC591, 16'hE564, 16'hF5A7, 16'h054E,
 16'h0DBD, 16'h1539, 16'h44D1, 16'h7825,
 16'h33E4, 16'hC714, 16'hB4F3, 16'hB807,
 16'hC5FE, 16'hE4FF, 16'hF002, 16'h00FF,
 16'h06FD, 16'h1009, 16'h43F1, 16'h6D16,
 16'h26E2, 16'hC326, 16'hB1D1, 16'hB73A,
 16'hCBBA, 16'hE651, 16'hF4A4, 16'h0566,
 16'h0B91, 16'h1578, 16'h447F, 16'h7089,
 16'h2970, 16'hC696, 16'hB765, 16'hBC9F,
 16'hD05F, 16'hE6A1, 16'hF361, 16'h039D,
 16'h0D65, 16'h0E99, 16'h3D68, 16'h6F96,
 16'h3A6E, 16'hD78E, 16'hB377, 16'hB983,
 16'hC682, 16'hE37A, 16'hF48A, 16'h0472,
 16'h0D92, 16'h0E6B, 16'h2C96, 16'h646B,
 16'h5393, 16'hF76F, 16'hBB90, 16'hB270,
 16'hC290, 16'hDB71, 16'hF18D, 16'hFE75,
 16'h0689, 16'h0C79, 16'h1B86, 16'h467B,
 16'h6E83, 16'h287F, 16'hC680, 16'hB781,
 16'hB980, 16'hCF7D, 16'hE986, 16'hF777,
 16'h048D, 16'h0A6F, 16'h0E95, 16'h2766,
 16'h5F9F, 16'h595C, 16'h03A9, 16'hBB53,
 16'hAEB1, 16'hC34B, 16'hD9B9, 16'hF042,
 16'hFCC4, 16'h0537, 16'h0ECC, 16'h1231,
 16'h2FD2, 16'h672B, 16'h4BD8, 16'hEB25,
 16'hB5DE, 16'hB320, 16'hC5E1, 16'hDE1D,
 16'hF0E6, 16'hFD18, 16'h0AEA, 16'h1014,
 16'h0FED, 16'h3511, 16'h67F3, 16'h4309,
 16'hE5FA, 16'hB903, 16'hB400, 16'hC6FD,
 16'hDF06, 16'hEEF6, 16'h010F, 16'h0AED,
 16'h0C16, 16'h0DE6, 16'h2E1E, 16'h60DF,
 16'h4C25, 16'hF1D6, 16'hB92E, 16'hB2CF,
 16'hC633, 16'hDDCC, 16'hEF34, 16'hFCCD,
 16'h0732, 16'h0DCE, 16'h0F31, 16'h23D2,
 16'h502B, 16'h5FD9, 16'h1122, 16'hBFE2,
 16'hB31A, 16'hBAEB, 16'hCF0F, 16'hEAF7,
 16'hFB03, 16'h0404, 16'h0BF5, 16'h0B11,
 16'h15E8, 16'h371F, 16'h64DB, 16'h3A2B,
 16'hD8CF, 16'hB636, 16'hB4C6, 16'hC83D,
 16'hDFC0, 16'hF342, 16'h00BD, 16'h0A43,
 16'h08BF, 16'h0D3E, 16'h1FC4, 16'h4539,
 16'h64CC, 16'h1B2F, 16'hC3D7, 16'hB321,
 16'hB5E7, 16'hCE10, 16'hE8FA, 16'hF5FC,
 16'h020E, 16'h06E8, 16'h0C21, 16'h10D7,
 16'h2130, 16'h4BC9, 16'h5C3F, 16'h14B9,
 16'hBF4E, 16'hB2AD, 16'hBE57, 16'hCEA5,
 16'hE85E, 16'hF7A0, 16'h0062, 16'h0B9E,
 16'h0D60, 16'h0AA1, 16'h205F, 16'h48A2,
 16'h5D5D, 16'h1BA5, 16'hBF58, 16'hB4AB,
 16'hBB52, 16'hCAB1, 16'hE64D, 16'hF6B5,
 16'h0249, 16'h0AB8, 16'h1047, 16'h0EBA,
 16'h1A46, 16'h3AB9, 16'h6049, 16'h30B5,
 16'hD94E, 16'hB5AF, 16'hB652, 16'hC5AE,
 16'hDE53, 16'hF3AC, 16'hFC55, 16'h08A9,
 16'h0E58, 16'h0DA9, 16'h0D55, 16'h23AE,
 16'h4B4E, 16'h57B7, 16'h0F43, 16'hBEC5,
 16'hB331, 16'hBDD9, 16'hD41D, 16'hE4EE,
 16'hF608, 16'h0201, 16'h06F5, 16'h0C16,
 16'h0DDE, 16'h132F, 16'h2AC4, 16'h5549,
 16'h45AB, 16'hF960, 16'hBB95, 16'hAF75,
 16'hC083, 16'hD785, 16'hEF75, 16'hF68E,
 16'h026F, 16'h0B94, 16'h096B, 16'h0B95,
 16'h0E6C, 16'h2791, 16'h5074, 16'h4986,
 16'hFF80, 16'hBC79, 16'hB090, 16'hC167,
 16'hD5A3, 16'hE952, 16'hF6B9, 16'h043D,
 16'h0ACC, 16'h0A2D, 16'h0ED9, 16'h0E21,
 16'h1FE5, 16'h4515, 16'h53F1, 16'h1709,
 16'hC5FC, 16'hB501, 16'hBC01, 16'hCDFE,
 16'hE500, 16'hF503, 16'h01FA, 16'h090B,
 16'h07EF, 16'h0916, 16'h0CE4, 16'h1223,
 16'h2CD6, 16'h5031, 16'h40C7, 16'hF442,
 16'hB7B5, 16'hB354, 16'hC6A3, 16'hD865,
 16'hEE94, 16'hFA72, 16'hFF89, 16'h087B,
 16'h0B82, 16'h0F81, 16'h117C, 16'h1287,
 16'h3076, 16'h538C, 16'h3773, 16'hEC8E,
 16'hB873, 16'hB28B, 16'hC576, 16'hDC89,
 16'hED79, 16'hFB85, 16'h077E, 16'h087F,
 16'h0884, 16'h0E79, 16'h0E89, 16'h1275,
 16'h2A8D, 16'h4973, 16'h458C, 16'hFF75,
 16'hBC8A, 16'hB276, 16'hBE8B, 16'hD475,
 16'hEB8A, 16'hF878, 16'h0385, 16'h0A7E,
 16'h0B7F, 16'h0E84, 16'h0E78, 16'h0C8C,
 16'h1671, 16'h3890, 16'h4F70, 16'h228F,
 16'hD873, 16'hB58A, 16'hB57A, 16'hCA81,
 16'hDE85, 16'hF075, 16'hFF91, 16'h0368,
 16'h0BA0, 16'h0A58, 16'h0EB1, 16'h0D45,
 16'h0BC5, 16'h1D31, 16'h36D9, 16'h4D1E,
 16'h1DEA, 16'hD40E, 16'hB9F9, 16'hB402,
 16'hC802, 16'hE1FB, 16'hF307, 16'h00F7,
 16'h0A09, 16'h0EF9, 16'h0E04, 16'h1101,
 16'h0BF8, 16'h0810, 16'h12E7, 16'h3023,
 16'h47D3, 16'h3437, 16'hEEBF, 16'hB84B,
 16'hB2AB, 16'hC55F, 16'hDB98, 16'hEE6F,
 16'hFC8B, 16'h0379, 16'h0B86, 16'h0E79,
 16'h0E89, 16'h0E72, 16'h0A96, 16'h0B60,
 16'h19AD, 16'h3644, 16'h4CCB, 16'h1C25,
 16'hD3EC, 16'hB602, 16'hB211, 16'hC5DC,
 16'hDB38, 16'hE9B3, 16'hFC61, 16'h048C,
 16'h0786, 16'h0D6B, 16'h0BA2, 16'h0852,
 16'h07B7, 16'h0644, 16'h0FBE, 16'h3342,
 16'h47BC, 16'h2248, 16'hE2B3, 16'hB654,
 16'hB1A1, 16'hCA6D, 16'hD984, 16'hEE8D,
 16'hFD61, 16'h03B0, 16'h0B3F, 16'h0AD2,
 16'h0F1E, 16'h0BF2, 16'h09FE, 16'h0911,
 16'h06E2, 16'h1C29, 16'h3BCF, 16'h4237,
 16'h0FC5, 16'hCB3D, 16'hB5C2, 16'hB73E,
 16'hCFC6, 16'hE333, 16'hF1D4, 16'h0424,
 16'h08E5, 16'h0E12, 16'h0DF8, 16'h0CFD,
 16'h0B0E, 16'h0BE7, 16'h0823, 16'h06D4,
 16'h1934, 16'h36C6, 16'h453F, 16'h18BD,
 16'hD445, 16'hB8BA, 16'hB746, 16'hCCBC,
 16'hE141, 16'hF2C3, 16'hFF38, 16'h08CE,
 16'h0E2B, 16'h0ADC, 16'h101C, 16'h09ED,
 16'h080A, 16'h08FE, 16'h0AFB, 16'h0E0C,
 16'h20EE, 16'h3917, 16'h37E4, 16'h0B20,
 16'hC8DE, 16'hB624, 16'hBEDB, 16'hCF24,
 16'hE4DF, 16'hF41B, 16'hFFED, 16'h0B0B,
 16'h0AFD, 16'h0AFA, 16'h100F, 16'h0AE8,
 16'h0B22, 16'h07D4, 16'h0635, 16'h07C3,
 16'h1544, 16'h2FB5, 16'h4052, 16'h20A7,
 16'hDF60, 16'hB99B, 16'hB467, 16'hCC98,
 16'hE068, 16'hF199, 16'hFB66, 16'h029C,
 16'h0E60, 16'h0AA6, 16'h0B52, 16'h0DB7,
 16'h0D3F, 16'h06CC, 16'h0929, 16'h06E2,
 16'h0111, 16'h15FD, 16'h2FF5, 16'h3C18,
 16'h1EDC, 16'hE42F, 16'hB9C6, 16'hB546,
 16'hC7AE, 16'hDB5C, 16'hED9D, 16'hFA69,
 16'h0591, 16'h0975, 16'h0D86, 16'h0E7E,
 16'h0D7F, 16'h0A83, 16'h077C, 16'h0884,
 16'h057E, 16'h027E, 16'h0386, 16'h1977,
 16'h2E8C, 16'h3870, 16'h1495, 16'hD666,
 16'hBC9E, 16'hB65F, 16'hCCA3, 16'hDE5B,
 16'hEFA8, 16'h0054, 16'h06B0, 16'h0A4D,
 16'h09B5, 16'h0E4A, 16'h0AB6, 16'h0B4B,
 16'h07B4, 16'h094C, 16'h06B4, 16'h044C,
 16'hFEB4, 16'h094E, 16'h20AE, 16'h3155,
 16'h36A8, 16'h035C, 16'hCAA1, 16'hB462,
 16'hBB9A, 16'hD06A, 16'hE492, 16'hF573,
 16'h0187, 16'h0780, 16'h0B79, 16'h0A8E,
 16'h0E6A, 16'h0B9F, 16'h0657, 16'h08B4,
 16'h0741, 16'h02C9, 16'hFF2E, 16'h04DC,
 16'hFE19, 16'h0CF2, 16'h2602, 16'h350A,
 16'h25EB, 16'hF320, 16'hC4D6, 16'hB631,
 16'hC1C9, 16'hD53C, 16'hEAC1, 16'hF741,
 16'h06BD, 16'h0843, 16'h0CC0, 16'h0E3C,
 16'h09CA, 16'h0E2D, 16'h0ADE, 16'h0416,
 16'h05F7, 16'h04FC, 16'h0111, 16'h01E2,
 16'hFD2B, 16'h00C7, 16'h1149, 16'h28A6,
 16'h356B, 16'h1C85, 16'hE889, 16'hC46B,
 16'hB7A0, 16'hC156, 16'hDAB3, 16'hEA46,
 16'hFABE, 16'h0440, 16'h07C1, 16'h0D3F,
 16'h0BC1, 16'h0B40, 16'h08BE, 16'h0A45,
 16'h04B8, 16'h004C, 16'h04AF, 16'h0256,
 16'hFCA5, 16'h0160, 16'h019D, 16'hFD65,
 16'h1199, 16'h2669, 16'h2F95, 16'h1F6C,
 16'hF095, 16'hC668, 16'hB69D, 16'hC05E,
 16'hD6A8, 16'hE850, 16'hF6B9, 16'h043E,
 16'h0ACB, 16'h0C2D, 16'h0BDA, 16'h081F,
 16'h0BE9, 16'h0A0D, 16'h01FD, 16'h03F9,
 16'h0110, 16'h00E9, 16'h031C, 16'h03E0,
 16'h0023, 16'hFDDA, 16'h0129, 16'h0AD5,
 16'h192C, 16'h26D5, 16'h2D29, 16'h0DDA,
 16'hDE22, 16'hC2E3, 16'hB918, 16'hC7EE,
 16'hDF0B, 16'hEEFD, 16'hFCFB, 16'h040C,
 16'h0AED, 16'h0E19, 16'h0AE2, 16'h0C24,
 16'h0AD4, 16'h0834, 16'h07C5, 16'h0242,
 16'h05B7, 16'h044E, 16'hFEAD, 16'h0059,
 16'hFEA2, 16'hFE63, 16'h0197, 16'hFD6F,
 16'h038B, 16'h167A, 16'h2182, 16'h2D82,
 16'h1F7C, 16'hF685, 16'hCE79, 16'hBB89,
 16'hC276, 16'hD38C, 16'hE573, 16'hF78D,
 16'h0073, 16'h068C, 16'h0B77, 16'h0B85,
 16'h0D80, 16'h0D7B, 16'h0B8A, 16'h0371,
 16'h0694, 16'h0166, 16'h01A0, 16'h045B,
 16'h00AB, 16'hFF4E, 16'hFDBA, 16'h023D,
 16'h00CC, 16'hFE2C, 16'hFBDC, 16'h021C,
 16'h08EC, 16'h1B0C, 16'h22FC, 16'h28FB,
 16'h120D, 16'hE4EC, 16'hCA1B, 16'hB9DF,
 16'hC826, 16'hD7D4, 16'hED32, 16'hF8C9,
 16'h023B, 16'h09C3, 16'h0C3E, 16'h0BC2,
 16'h0A3D, 16'h08C5, 16'h0738, 16'h08CC,
 16'h012F, 16'h06D7, 16'h0322, 16'hFFE6,
 16'h0111, 16'hFFF9, 16'h03FC, 16'h0010,
 16'hFDE3, 16'hFF2A, 16'hFCCA, 16'h0141,
 16'h01B4, 16'hFF58, 16'h069B, 16'h1571,
 16'h1E84, 16'h2385, 16'h2275, 16'hFD8F,
 16'hD96F, 16'hC191, 16'hBD70, 16'hCB8E,
 16'hDD77, 16'hF381, 16'hFA88, 16'h046E,
 16'h0A9E, 16'h0E55, 16'h0DB9, 16'h0C37,
 16'h0ADB, 16'h0112, 16'h0401, 16'hFFEC,
 16'h0027, 16'hFFC6, 16'hFA4D, 16'h00A1,
 16'h006F, 16'hFC83, 16'hFA89, 16'hFD6D,
 16'hFE9B, 16'hFC5E, 16'hFDA8, 16'h0055,
 16'hFCAB, 16'hFC58, 16'hFCA2, 16'hFD66,
 16'h0691, 16'h0E79, 16'h197C, 16'h1E91,
 16'h1C5F, 16'h06B2, 16'hE53D, 16'hCDD4,
 16'hBC1A, 16'hC6F9, 16'hD8F3, 16'hE921,
 16'hF7CB, 16'h0048, 16'h08A7, 16'h0A69,
 16'h0E88, 16'h0D84, 16'h0D73, 16'h0B95,
 16'h0A64, 16'h08A2, 16'h0259, 16'h00AA,
 16'h0357, 16'h00A5, 16'hFE61, 16'h0498,
 16'hFE70, 16'hFE87, 16'h0384, 16'hFD70,
 16'hFD9C, 16'h0158, 16'hFFB3, 16'hFD43,
 16'hFDC7, 16'hFE2F, 16'hFFDA, 16'h001E,
 16'hFFE9, 16'hFD12, 16'h00F2, 16'h020A,
 16'h0AF8, 16'h1808, 16'h17F6, 16'h1C0E,
 16'h15ED, 16'hFE19, 16'hE2E0, 16'hD228,
 16'hC0CE, 16'hC53C, 16'hD8BB, 16'hE94D,
 16'hF7AC, 16'h045B, 16'h0A9E, 16'h0C68,
 16'h0E92, 16'h0C73, 16'h0A8A, 16'h0977,
 16'h098A, 16'h0473, 16'h0791, 16'h046B,
 16'h009A, 16'hFF5F, 16'h04A9, 16'h014E,
 16'hFFBD, 16'h0338, 16'hFFD2, 16'hFD24,
 16'hFCE5, 16'h0113, 16'hFEF4, 16'h0406,
 16'hFF00, 16'hFDF9, 16'h010D, 16'hFDEF,
 16'hFD14, 16'hFDEB, 16'hFC14, 16'hFCED,
 16'hFC13, 16'hFDEE, 16'h0010, 16'hFFF3,
 16'h0008, 16'hFFFE, 16'hFFFC, 16'h000A,
 16'h0DF1, 16'h0F13, 16'h14E9, 16'h131A,
 16'h0EE4, 16'h051E, 16'hEAE1, 16'hDB20,
 16'hCDDF, 16'hC621, 16'hCCE0, 16'hE01D,
 16'hE9E7, 16'hFB15, 16'h04EF, 16'h0B0D,
 16'h0FF6, 16'h0B06, 16'h0C00, 16'h09FA,
 16'h090B, 16'h0AF0, 16'h0314, 16'h18EA,
 16'h2F18, 16'hF6E6, 16'hE51B, 16'hF0E5,
 16'hF01A, 16'hF3E8, 16'h0115, 16'h25EF,
 16'hFA0C, 16'hE1FA, 16'h01FE, 16'hF00B,
 16'h03EB, 16'h2621, 16'hF5D3, 16'hE639,
 16'h01BA, 16'hEE53, 16'h07A1, 16'h256B,
 16'hF28B, 16'hE87E, 16'h007A, 16'hEF8C,
 16'h026F, 16'h2094, 16'hF76C, 16'hE592,
 16'hFF72, 16'hF388, 16'h007F, 16'h2078,
 16'hF694, 16'hE55E, 16'hFFB3, 16'hED39,
 16'h00DC, 16'h230E, 16'hF70B, 16'hE7DB,
 16'h0040, 16'hEBA4, 16'h0277, 16'h236F,
 16'hF3AB, 16'hE43C, 16'h00DC, 16'hEE0E,
 16'h0205, 16'h22EA, 16'hF425, 16'hEACF,
 16'h013A, 16'hEDBF, 16'h0046, 16'h1DB8,
 16'hF747, 16'hEEBC, 16'h013F, 16'hEDC9,
 16'hFD2C, 16'h1BE0, 16'hF911, 16'hF302,
 16'hFFEA, 16'hE92A, 16'hFDC1, 16'h1554,
 16'h0297, 16'hFA7F, 16'hF86A, 16'hEEAD,
 16'hF83D, 16'h0AD8, 16'h1214, 16'hFDFF,
 16'hF0EE, 16'hF324, 16'hF6CC, 16'h0442,
 16'h18B1, 16'hFE5A, 16'hE89C, 16'hF86D,
 16'hEF8B, 16'h047C, 16'h1E7E, 16'hFA86,
 16'hE477, 16'h008A, 16'hEB78, 16'hFE85,
 16'h227F, 16'hF37B, 16'hED8C, 16'h016B,
 16'hEC9F, 16'hFD57, 16'h19B4, 16'hFC41,
 16'hF6C9, 16'hFA2D, 16'hEEDE, 16'hF717,
 16'h0AF4, 16'h1101, 16'hFE0A, 16'hECED,
 16'hF71A, 16'hF3E0, 16'h0425, 16'h22D8,
 16'hF629, 16'hE4D7, 16'h0027, 16'hEBDE,
 16'hFD1C, 16'h22EA, 16'hF60E, 16'hEBFB,
 16'hFFFB, 16'hEE11, 16'hFCE3, 16'h1428,
 16'h01CD, 16'hFA3E, 16'hF5B7, 16'hF354,
 16'hF9A2, 16'h0367, 16'h1E92, 16'h0073,
 16'hEA8A, 16'hFD76, 16'hED8D, 16'h046F,
 16'h2396, 16'hF564, 16'hECA3, 16'h0154,
 16'hEDB7, 16'hFD3D, 16'h15CF, 16'h0325,
 16'hFFE7, 16'hF60D, 16'hEFFE, 16'hF5F9,
 16'h040F, 16'h1DEA, 16'hFB1B, 16'hE8E1,
 16'h0022, 16'hEEDD, 16'h0022, 16'h1EE1,
 16'hF719, 16'hF5EF, 16'hFC08, 16'hF001,
 16'hF9F7, 16'h0A12, 16'h15E3, 16'hFE28,
 16'hEDCD, 16'hFD3E, 16'hF1B9, 16'h014E,
 16'h22AC, 16'hF459, 16'hEFA3, 16'hFF5F,
 16'hEEA2, 16'hFC5B, 16'h0FAA, 16'h0D4F,
 16'hFFB9, 16'hF03E, 16'hF5CD, 16'hF326,
 16'h01E9, 16'h2306, 16'hF80C, 16'hE9E2,
 16'hFD30, 16'hF2BF, 16'hFD51, 16'h11A0,
 16'h0A6F, 16'hFA82, 16'hF08C, 16'hF968,
 16'hF3A2, 16'h0156, 16'h25AF, 16'hF54E,
 16'hE9B4, 16'h004C, 16'hF0B1, 16'hFB53,
 16'h10A8, 16'h0D5F, 16'h0199, 16'hF370,
 16'hF685, 16'hF588, 16'h016A, 16'h1FA4,
 16'hF34E, 16'hF3BF, 16'hFD35, 16'hF2D7,
 16'hFE1E, 16'h03EB, 16'h1A0C, 16'hFEFD,
 16'hECFC, 16'hFD09, 16'hF3F2, 16'hFF12,
 16'h18EB, 16'hFD18, 16'hF7E6, 16'hF71A,
 16'hF5E7, 16'hF716, 16'h03ED, 16'h2610,
 16'hF8F5, 16'hED06, 16'hFCFD, 16'hF000,
 16'hF702, 16'h07FE, 16'h0B02, 16'hFBFE,
 16'hED01, 16'hF301, 16'hF4FD, 16'hFB07,
 16'h18F3, 16'hFA13, 16'hF3E7, 16'hF721,
 16'hEFD6, 16'hF933, 16'h00C3, 16'h2247,
 16'hF6B1, 16'hEB56, 16'hFAA3, 16'hF063,
 16'hFB99, 16'h0869, 16'h1697, 16'hFE67,
 16'hEF9D, 16'hFA5E, 16'hF4A8, 16'hFA50,
 16'h14BA, 16'h0439, 16'hFBD8, 16'hF715,
 16'hF2FF, 16'hF3EB, 16'h022B, 16'h1BC1,
 16'hF754, 16'hF596, 16'hFA80, 16'hF56A,
 16'hF9AB, 16'h0343, 16'h1FCD, 16'hF725,
 16'hECE7, 16'hFC0F, 16'hF2F8, 16'hFC04,
 16'h08FF, 16'h1B00, 16'hFAFD, 16'hEE0A,
 16'hFAEC, 16'hF521, 16'hFDD1, 16'h0A3E,
 16'h0DB1, 16'hFF61, 16'hF38B, 16'hF68B,
 16'hF55F, 16'hFFB8, 16'h1230, 16'h03E7,
 16'hF904, 16'hF310, 16'hF5DE, 16'hFA31,
 16'hFFC3, 16'h1748, 16'hFFAF, 16'hF757,
 16'hFCA4, 16'hF360, 16'hF39F, 16'h0360,
 16'h18A2, 16'hF75A, 16'hF7AD, 16'hFA4A,
 16'hF5C0, 16'hF936, 16'hFFD5, 16'h1C1F,
 16'hF9ED, 16'hF708, 16'hFC02, 16'hF6F4,
 16'hFA16, 16'h00E0, 16'h1E29, 16'hF3CF,
 16'hF337, 16'hFDC5, 16'hF63E, 16'hFAC0,
 16'h0041, 16'h1EBF, 16'hF440, 16'hF2C2,
 16'hFE3C, 16'hF6C7, 16'hF734, 16'h03D3,
 16'h1E26, 16'hF3E0, 16'hF61A, 16'hFCEA,
 16'hF614, 16'hF7ED, 16'h0412, 16'h19EE,
 16'hF612, 16'hF5EE, 16'hFA13, 16'hF9EB,
 16'hFB18, 16'hFFE3, 16'h1924, 16'hF6D4,
 16'hF835, 16'hFAC3, 16'hF544, 16'hF9B5,
 16'h0052, 16'h16A7, 16'hF860, 16'hFC99,
 16'hFC6D, 16'hF38E, 16'hFA76, 16'hFD88,
 16'h1078, 16'h0089, 16'hF875, 16'hF68F,
 16'hF16C, 16'hF899, 16'hFE62, 16'h0EA5,
 16'h0952, 16'hF9B8, 16'hF53C, 16'hF5D1,
 16'hFB23, 16'hF6E9, 16'h070A, 16'h1204,
 16'hFCEC, 16'hF725, 16'hF6CB, 16'hF945,
 16'hF7AC, 16'h0361, 16'h1992, 16'hF97B,
 16'hF27A, 16'hFA90, 16'hF566, 16'hF7A3,
 16'h0256, 16'h1AAF, 16'hF54E, 16'hF1B3,
 16'hFA4D, 16'hF2B4, 16'hFD4B, 16'h03B5,
 16'h114C, 16'hF9B2, 16'hFC52, 16'hFAAA,
 16'hF15A, 16'hFAA0, 16'hFB67, 16'h0992,
 16'h0D76, 16'hFE83, 16'hF682, 16'hF679,
 16'hFC8B, 16'hF773, 16'h038F, 16'h1A70,
 16'hF890, 16'hF371, 16'hFC8C, 16'hFB78,
 16'hF883, 16'h0183, 16'h1777, 16'hFA8F,
 16'hF56A, 16'hFD9D, 16'hF65B, 16'hFAAD,
 16'hFD4B, 16'h0ABD, 16'h0D3C, 16'hFACA,
 16'hF632, 16'hF6CF, 16'hFC32, 16'hF5CC,
 16'h0338, 16'h19C3, 16'hF544, 16'hF5B2,
 16'hFC5A, 16'hF398, 16'hFD7A, 16'hFE72,
 16'h0AA3, 16'h0446, 16'hFBD2, 16'hFB16,
 16'hF404, 16'hFAE1, 16'hF738, 16'h03B1,
 16'h1A65, 16'hF887, 16'hF18D, 16'hF860,
 16'hF6B0, 16'hF843, 16'hFFC7, 16'h1132,
 16'hFDD4, 16'hFA28, 16'hF9D9, 16'hF229,
 16'hFDD1, 16'hF738, 16'h03BC, 16'h1853,
 16'hF39D, 16'hF374, 16'hFA7A, 16'hF596,
 16'hF95B, 16'hFFB4, 16'h0E3F, 16'hFFCC,
 16'hFB29, 16'hFBE0, 16'hF41B, 16'hF9E8,
 16'hF817, 16'h02E7, 16'h191E, 16'hF3DB,
 16'hF42F, 16'hFFC4, 16'hF44B, 16'hFDA6,
 16'hFD6A, 16'h0A83, 16'h0891, 16'hF95A,
 16'hF7BD, 16'hF62C, 16'hF9E9, 16'hF703,
 16'h040F, 16'h13E2, 16'hF82B, 16'hFBCA,
 16'hFD3D, 16'hF2BE, 16'h0145, 16'hF8BB,
 16'h0143, 16'h17C1, 16'hFB37, 16'hF5D5,
 16'hFD1C, 16'hF5F5, 16'hFFF9, 16'hFA1A,
 16'h08D1, 16'h0F47, 16'hFF9E, 16'hF77E,
 16'hF566, 16'hF9B6, 16'hFB2E, 16'hFFEE,
 16'h0DF6, 16'hFE26, 16'hF8C0, 16'hFD59,
 16'hF58F, 16'h0188, 16'hF461, 16'h04B5,
 16'h1337, 16'hF7DB, 16'hF916, 16'hFDF6,
 16'hF600, 16'h0109, 16'hF8EF, 16'h0117,
 16'h17E5, 16'hF91D, 16'hF6E4, 16'hFE19,
 16'hF4EC, 16'h020C, 16'hFDFD, 16'h01F9,
 16'h1412, 16'hFAE4, 16'hF826, 16'hFDCE,
 16'hF63F, 16'h01B4, 16'hFB59, 16'h049B,
 16'h0971, 16'hFA83, 16'hF788, 16'hF76E,
 16'hFC9B, 16'hFD5E, 16'h00A8, 16'h0C52,
 16'h08B5, 16'h0045, 16'hF7BF, 16'hF83D,
 16'hFDC7, 16'hFE37, 16'hFDCB, 16'h0832,
 16'h08D0, 16'hFA2F, 16'hF9D3, 16'hFC2B,
 16'hFCD7, 16'hFD26, 16'h00DE, 16'h061D,
 16'h08E8, 16'hFF14, 16'hF7F0, 16'hF70C,
 16'hFAF8, 16'h0003, 16'h0002, 16'h06FA,
 16'h090A, 16'hFCF2, 16'hF811, 16'hFBEC,
 16'hFC17, 16'hFCE6, 16'hFC1C, 16'h06E3,
 16'h0C1C, 16'hFEE7, 16'hF815, 16'hFCF0,
 16'hFC0A, 16'hFCFC, 16'hFCFE, 16'h0409,
 16'h0FF0, 16'hFF17, 16'hF2E1, 16'hF727,
 16'hF2D1, 16'hFA37, 16'hFAC2, 16'h0044,
 16'h0FB6, 16'hF54F, 16'hF2AE, 16'hFC54,
 16'hF5AB, 16'hFE53, 16'hF6B1, 16'h024A,
 16'h0FBD, 16'hF53A, 16'hF9D0, 16'h0025,
 16'hF2E8, 16'h0009, 16'hF908, 16'h00E5,
 16'h0B31, 16'hF7B7, 16'hFD62, 16'hFC85,
 16'hF695, 16'hFF51, 16'hFBC9, 16'h001D,
 16'h07FC, 16'h02EE, 16'hFD27, 16'hFBC4,
 16'hFB4E, 16'hF8A2, 16'h016C, 16'hFD89,
 16'h027F, 16'h0C7B, 16'hFC88, 16'hF779,
 16'hFE81, 16'hF989, 16'h006C, 16'hFBA1,
 16'hFD4F, 16'h0CC3, 16'hF828, 16'hFBF0,
 16'hFCF7, 16'hFA22, 16'hFFC3, 16'hFF58,
 16'h008D, 16'h038E, 16'h0759, 16'hFDBD,
 16'hF92F, 16'hFCE4, 16'hFA0B, 16'h0003,
 16'hFBF2, 16'h0116, 16'h0EE6, 16'hF61B,
 16'hFBE5, 16'hFD19, 16'hF9EB, 16'h0010,
 16'hFFF6, 16'h0002, 16'h0307, 16'h07EF,
 16'hFD1A, 16'hF8DF, 16'hFD27, 16'hF9D4,
 16'h0030, 16'hFECC, 16'h0137, 16'h0DC8,
 16'hF739, 16'hFCC7, 16'hFC37, 16'hFACD,
 16'hFF2D, 16'hFFDA, 16'hFF1F, 16'h00E9,
 16'h080F, 16'hFDF8, 16'hFA01, 16'hFC05,
 16'hFCF6, 16'hFC0F, 16'hFDEE, 16'h0112,
 16'h0CF0, 16'hFA0B, 16'hFCFC, 16'hFCFD,
 16'hFA0B, 16'hFFEB, 16'hFD21, 16'hFED0,
 16'h0141, 16'h0CAF, 16'hF761, 16'hF98E,
 16'hFD82, 16'hFA6F, 16'hFBA1, 16'hFF51,
 16'hFFBA, 16'h003C, 16'h08CC, 16'hFC2E,
 16'hFCD6, 16'hFC29, 16'hFAD6, 16'hFF2D,
 16'hFFCD, 16'hFF3B, 16'h04BC, 16'h014E,
 16'hFAA7, 16'hFC65, 16'hFC8E, 16'hFC80,
 16'hFD71, 16'hFD9E, 16'hFD54, 16'h07B9,
 16'hFD3A, 16'hFCD1, 16'hFC26, 16'hFAE2,
 16'hFB17, 16'hFEEE, 16'h000F, 16'hFEF1,
 16'h0912, 16'hF6E9, 16'hFB1D, 16'hF9DD,
 16'hFB29, 16'hFCD0, 16'h0039, 16'hFFBD,
 16'hFF4E, 16'h08A7, 16'hF863, 16'hFB93,
 16'hFD76, 16'hFB83, 16'hFB84, 16'hFF77,
 16'hFF8A, 16'hFF77, 16'h0787, 16'hFA7D,
 16'hFA7E, 16'hFF86, 16'hF677, 16'hFC8D,
 16'h006E, 16'hFE98, 16'h005F, 16'h06AC,
 16'hFB4A, 16'hF9C0, 16'h0036, 16'hF9D3,
 16'hFB25, 16'hFAE2, 16'hFA19, 16'h00EB,
 16'h0811, 16'hF9F2, 16'hFD0C, 16'hFBF4,
 16'hF70E, 16'hFFEF, 16'h0015, 16'hF9E5,
 16'h0220, 16'h06DB, 16'h012B, 16'h01CF,
 16'hF836, 16'hFBC5, 16'hFD40, 16'hFBBA,
 16'hFD4D, 16'hFBAC, 16'h015B, 16'h05A0,
 16'hFD63, 16'hFC9A, 16'hFD69, 16'hFC94,
 16'hFA6E, 16'hFF92, 16'hFF6E, 16'hFF91,
 16'h086F, 16'hF792, 16'hFA6D, 16'hFF95,
 16'hFC69, 16'hFF99, 16'h0064, 16'hFBA1,
 16'hFD59, 16'h02AE, 16'hFD4A, 16'hFBBD,
 16'hFD3D, 16'hFCC9, 16'hFD31, 16'hFDD5,
 16'hFE23, 16'hFCE6, 16'hFE11, 16'h07F8,
 16'hFCFF, 16'hF80A, 16'hFCEC, 16'hFD1F,
 16'hFAD5, 16'hFF37, 16'hFFBF, 16'hFF48,
 16'h07B2, 16'hFA54, 16'hFCA7, 16'hFC5D,
 16'hFAA1, 16'hFF5E, 16'hFAA5, 16'h0057,
 16'hFEAF, 16'h004A, 16'h03BF, 16'hFE35,
 16'hFBD9, 16'hFD18, 16'hFBF9, 16'hFAF5,
 16'hFF1D, 16'hFAD1, 16'hFF42, 16'h04AB,
 16'hFA67, 16'hFC87, 16'hFD8A, 16'hF967,
 16'h00A8, 16'hFF4A, 16'hFFC2, 16'hFF32,
 16'h00D9, 16'h061F, 16'hFAE7, 16'hFC15,
 16'hFCED, 16'hFC12, 16'hFCED, 16'hFD16,
 16'hFDE5, 16'hFD21, 16'h02D9, 16'h052E,
 16'hFDC8, 16'hFB44, 16'hFDAE, 16'hFB61,
 16'hFD91, 16'hFC7C, 16'hFE76, 16'hFD99,
 16'h0159, 16'h01B4, 16'hFC3F, 16'hFCCE,
 16'hFC25, 16'hFCE9, 16'hFD09, 16'hFE04,
 16'hFCEF, 16'hFE1D, 16'h00D8, 16'h0133,
 16'hFBC4, 16'hFD42, 16'hFCB9, 16'hFC4B,
 16'hFDB3, 16'hFD4F, 16'hFDAF, 16'hFD51,
 16'h03B1, 16'hFD4C, 16'hFBB9, 16'hFD41,
 16'hFBC5, 16'hFE33, 16'hFCD6, 16'hFE21,
 16'hFCEA, 16'h0209, 16'h0104, 16'hFAEE,
 16'h0021, 16'hFCD2, 16'hFC3A, 16'h00BA,
 16'hFC52, 16'hFCA2, 16'hFC6A, 16'hFC8C,
 16'h017C, 16'hFF7D, 16'hFD89, 16'hFC72,
 16'hFC92, 16'hFC6D, 16'hFD90, 16'hFD75,
 16'hFD84, 16'h0185, 16'h0172, 16'h0198,
 16'hFD5C, 16'hFCB1, 16'hFC40, 16'hFCD1,
 16'hFD1D, 16'hFCF5, 16'h00F9, 16'hFC1A,
 16'h00D2, 16'h0641, 16'hFCAC, 16'hFD66,
 16'h008B, 16'hFD82, 16'hFC71, 16'hFC9B,
 16'h005B, 16'hFCAD, 16'h004D, 16'h02B8,
 16'hF945, 16'hFDBB, 16'hFF47, 16'hFDB5,
 16'hFF52, 16'hFDA6, 16'hFB62, 16'hFD94,
 16'h0077, 16'h007E, 16'h018D, 16'hFA68,
 16'hFCA2, 16'hFC53, 16'hFCB8, 16'hFD3E,
 16'hFDCB, 16'hFE2D, 16'hF8DA, 16'h0120,
 16'hFFE4, 16'hFA1A, 16'hFAE7, 16'hFA1A,
 16'hF9E4, 16'hFD1E, 16'hF9DD, 16'hFE2B,
 16'hFECC, 16'hFB3E, 16'hFEB7, 16'h0053,
 16'hFEA3, 16'hFB68, 16'hFE8D, 16'hFB7D,
 16'hFE7A, 16'h008E, 16'hFE6C, 16'h009A,
 16'hFE5F, 16'h01A7, 16'h0055, 16'hFCAD,
 16'h0053, 16'hFCAB, 16'hFC59, 16'hFCA2,
 16'hFC64, 16'hFE94, 16'hFC75, 16'hFE82,
 16'h0088, 16'hFD6D, 16'hFC9E, 16'hFC58,
 16'hFDB2, 16'hFE44, 16'hFDC5, 16'hFE33,
 16'hFED4, 16'h0026, 16'hFFE0, 16'h011A,
 16'hFCEB, 16'hFD11, 16'hFCF2, 16'hFC0C,
 16'hFDF4, 16'hFD0D, 16'hFDF1, 16'hFD12,
 16'hFDEB, 16'h0117, 16'h00E6, 16'hFD1E,
 16'hFBDE, 16'hFD25, 16'hFCD9, 16'h0129,
 16'hFCD5, 16'hFC2C, 16'h00D3, 16'hFC2E,
 16'h00D2, 16'h002D, 16'hFCD4, 16'hFD2C,
 16'hFCD4, 16'hFC2C, 16'hFDD4, 16'hFD2B,
 16'hFDD6, 16'h012A, 16'hFCD5, 16'hFC2D,
 16'h00CF, 16'hFC36, 16'hFCC5, 16'hFD40,
 16'hFBBA, 16'h024C, 16'hFBAF, 16'hFD57,
 16'hFBA2, 16'hFD65, 16'h0094, 16'hFD73,
 16'h0086, 16'hFD81, 16'h0078, 16'h018E,
 16'hFC6D, 16'hFD98, 16'hFF64, 16'hFD9E,
 16'hFF61, 16'hFDA0, 16'hFF61, 16'h019C,
 16'hFC68, 16'hFC93, 16'hFC74, 16'hFC84,
 16'h0085, 16'hFC70, 16'hFC9C, 16'hFC58,
 16'hFDB4, 16'hFF40, 16'hFFCC, 16'h0028,
 16'hFCE5, 16'h010D, 16'hFD01, 16'hFCF1

};

logic [17:0] shoot_depth;
logic shoot_repeats;
assign shoot_depth = 18'd4080; // same as numbers of samples
assign shoot_repeats = 1;
/* end sine 441 hz*/
assign dout[15:0] = shoot_ROM[adress][15:0];
assign repeats = shoot_repeats;
assign depth = shoot_depth;


endmodule 