module semi_ROM (
	
	input clk,
	input resetN,
	//input read, // current word is being read
	//input next_word // current word was done being read
	input [8:0] adress, // for future purpose
	output [15:0] dout,
	output [17:0] depth,
	output repeats

);
/*sawing pattern
wire [9:0][15:0] ROM; // stroe the value
wire [15:0] counter; // 
wire rom_full;
assign depth = 10; // there are 10 rows (for now)

always_ff @(posedge clk, negedge resetN) begin
    if(resetN == 1'b0) begin
		//dout <= 0;
		//repeats <= 0;
		counter <= 16'b0;
		rom_full <= 0;
	 end
	 else begin
		 if (counter <= 16'd9 && rom_full == 0) begin // fill the Rom once
			counter <= counter + 1;
			ROM[counter][15:0] <= counter;
		 end
		 else begin
			rom_full <= 1;
		 end
	 end

end*/


///* sine 440 hz - one cycle*/
// // stroe the value
//logic [0:99][15:0] ROM ={ // need to be 0 to 102 so first 2 bytes be on the left 
// 16'h0380, 16'h09e8, 16'h1045, 16'h1694, 16'h1cc8, 16'h22e3, 16'h28d9, 16'h2ea6, 16'h3447, 16'h39ad, 16'h3ee2, 16'h43cb, 16'h4881, 16'h4cdc, 16'h50f9, 16'h54b9, 16'h582b, 16'h5b41, 16'h5dfe, 16'h6058, 16'h6257, 16'h63ec, 16'h6522, 16'h65f2, 16'h6658, 16'h665c, 16'h65f3, 16'h6528, 16'h63f5, 16'h6261, 16'h6065, 16'h5e0c, 16'h5b52, 16'h583d, 16'h54d1, 16'h510c, 16'h4cf8, 16'h4898, 16'h43ea, 16'h3efe, 16'h39cd, 16'h3466, 16'h2ec7, 16'h28fc, 16'h2306, 16'h1ced, 16'h16b7, 16'h106a, 16'h0a0c, 16'h03a8, 16'hfd38, 16'hf6d4, 16'hf072, 16'hea23, 16'he3ed, 16'hddc9, 16'hd7d7, 16'hd1fb, 16'hcc60, 16'hc6e8, 16'hc1b8, 16'hbcba, 16'hb80b, 16'hb399, 16'haf7f, 16'habad, 16'ha837, 16'ha512, 16'ha251, 16'h9fe2, 16'h9de4, 16'h9c39, 16'h9afd, 16'h9a22, 16'h99ac, 16'h99a2, 16'h99fb, 16'h9abb, 16'h9be3, 16'h9d6c, 16'h9f5d, 16'ha1ab, 16'ha459, 16'ha766, 16'haac6, 16'hae84, 16'hb28a, 16'hb6e9, 16'hbb87, 16'hc072, 16'hc597, 16'hcafb, 16'hd094, 16'hd656, 16'hdc4f, 16'he25c, 16'he897, 16'heeda, 16'hf53c, 16'hfb9d 
//
//};
//assign depth = 100; // same as numbers of row
///* end sine 440 hz*/



///* sine 440 hz - one second*/
// // stroe the value
//logic [0:705599] ROM =// need to be 0 to 102 so first 2 bytes be on the left 
//  
//;
//assign depth = 44100; // same as numbers of row
///* end sine 440 hz - one second*/




///* sine 441 hz - one cycle*/
// // stroe the value
//logic [0:98][15:0] ROM ={ // need to be 0 to 102 so first 2 bytes be on the left 
//16'h0000, 16'h066e, 16'h0cd6, 16'h132f,
// 16'h1979, 16'h1fa3, 16'h25b4, 16'h2b98,
// 16'h3156, 16'h36dd, 16'h3c32, 16'h4144,
// 16'h461c, 16'h4aa2, 16'h4ee9, 16'h52d6,
// 16'h5677, 16'h59bb, 16'h5ca9, 16'h5f33,
// 16'h6166, 16'h632c, 16'h6498, 16'h6598,
// 16'h6631, 16'h6668, 16'h6631, 16'h6599,
// 16'h6496, 16'h632e, 16'h6164, 16'h5f35,
// 16'h5ca8, 16'h59bc, 16'h5675, 16'h52d8,
// 16'h4ee6, 16'h4aa7, 16'h4617, 16'h4148,
// 16'h3c2e, 16'h36e0, 16'h3154, 16'h2b9a,
// 16'h25b2, 16'h1fa5, 16'h1977, 16'h1330,
// 16'h0cd6, 16'h066d, 16'h0001, 16'hf991,
// 16'hf32c, 16'heccf, 16'he688, 16'he05d,
// 16'hda4b, 16'hd46a, 16'hcea9, 16'hc922,
// 16'hc3cf, 16'hbebc, 16'hb9e5, 16'hb55d,
// 16'hb117, 16'had29, 16'ha98b, 16'ha644,
// 16'ha358, 16'ha0cb, 16'h9e9c, 16'h9cd2,
// 16'h9b69, 16'h9a69, 16'h99cd, 16'h999a,
// 16'h99cd, 16'h9a68, 16'h9b6a, 16'h9cd2,
// 16'h9e9b, 16'ha0cd, 16'ha356, 16'ha645,
// 16'ha98c, 16'had25, 16'hb11d, 16'hb558,
// 16'hb9e8, 16'hbeba, 16'hc3d1, 16'hc91f,
// 16'hceae, 16'hd463, 16'hda51, 16'he059,
// 16'he68c, 16'heccc, 16'hf32d
//
//};
//assign depth = 99; // same as numbers of samples
///* end sine 441 hz*/










///* sine 1000 hz*/
// // stroe the value
//logic [0:15][15:0] ROM ={ // need to be 0 to 102 so first 2 bytes be on the left 
//	16'h0f82, 16'h5009,
//	 16'h65b3, 16'h4337,
//	 16'hfa20, 16'hb559,
//	 16'h9927, 16'hb890,
//};
//assign depth = 16; // same as numbers of row
///* end sine 1000 hz*/


///* sine 1000 hz -  one second*/
// // stroe the value
//logic [0:44099][15:0] ROM ={ // need to be 0 to 102 so first 2 bytes be on the left 
//16'h2020, 16'h0e8a, 16'h1cca, 16'h2a72,
// 16'h3741, 16'h42ed, 16'h4d44, 16'h5602,
// 16'h5d0c, 16'h6229, 16'h6551, 16'h6664,
// 16'h656b, 16'h625f, 16'h5d57, 16'h5669,
// 16'h4dbd, 16'h437a, 16'h37df, 16'h2b1a,
// 16'h1d7f, 16'h0f41, 16'h20bb, 16'hf22f,
// 16'he3ea, 16'hd639, 16'hc95d, 16'hbd9e,
// 16'hb339, 16'haa62, 16'ha345, 16'h9e0c,
// 16'h9acb, 16'h999b, 16'h9a7e, 16'h9d6d,
// 16'ha25d, 16'ha933, 16'hb1cb, 16'hbbf7,
// 16'hc78a, 16'hd437, 16'he1d4, 16'hf002,
// 16'hfe8d, 16'h0d16, 16'h1b64, 16'h291c,
// 16'h3604, 16'h41d4, 16'h4c49, 16'h553a,
// 16'h5c69, 16'h61be, 16'h6518, 16'h6660,
// 16'h659e, 16'h62c1, 16'h5df1, 16'h572d,
// 16'h4eb0, 16'h4490, 16'h3917, 16'h2c6c,
// 16'h1ee2, 16'h10b4, 16'h0230, 16'hf3a1,
// 16'he553, 16'hd78c, 16'hca9c, 16'hbebd,
// 16'hb431, 16'hab33, 16'ha3e3, 16'h9e7d,
// 16'h9b06, 16'h99a3, 16'h9a4e, 16'h9d0b,
// 16'ha1c8, 16'ha870, 16'hb0da, 16'hbae5,
// 16'hc64f, 16'hd2ec, 16'he06b, 16'hee95,
// 16'hfd15, 16'h0ba6, 16'h19f8, 16'h27c8,
// 16'h34c5, 16'h40b1, 16'h4b53, 16'h5463,
// 16'h5bcb, 16'h6149, 16'h64da, 16'h6658,
// 16'h65c7, 16'h6326, 16'h5e7d, 16'h57f5,
// 16'h4f97, 16'h45a8, 16'h3a49, 16'h2dbd,
// 16'h2044, 16'h1225, 16'h03a4, 16'hf516,
// 16'he6ba, 16'hd8e6, 16'hcbdb, 16'hbfdf,
// 16'hb52f, 16'hac04, 16'ha48b, 16'h9ef0,
// 16'h9b48, 16'h99af, 16'h9a23, 16'h9cb0,
// 16'ha136, 16'ha7b2, 16'haff0, 16'hb9d1,
// 16'hc51e, 16'hd19c, 16'hdf0a, 16'hed25,
// 16'hfba1, 16'h0a2f, 16'h1893, 16'h266a,
// 16'h3387, 16'h3f8d, 16'h4a52, 16'h5391,
// 16'h5b1e, 16'h60d7, 16'h6493, 16'h664b,
// 16'h65ee, 16'h637f, 16'h5f0d, 16'h58af,
// 16'h5081, 16'h46ba, 16'h3b78, 16'h2f0c,
// 16'h21a4, 16'h1394, 16'h051b, 16'hf688,
// 16'he825, 16'hda41, 16'hcd1d, 16'hc104,
// 16'hb630, 16'hacdb, 16'ha537, 16'h9f68,
// 16'h9b8f, 16'h99bf, 16'h9a02, 16'h9c54,
// 16'ha0af, 16'ha6f3, 16'haf0c, 16'hb8c2,
// 16'hc3ee, 16'hd050, 16'hddaa, 16'hebb6,
// 16'hfa2b, 16'h08bc, 16'h1728, 16'h250d,
// 16'h3246, 16'h3e63, 16'h4953, 16'h52b4,
// 16'h5a73, 16'h605b, 16'h6448, 16'h663b,
// 16'h660b, 16'h63d7, 16'h5f96, 16'h5965,
// 16'h5169, 16'h47c2, 16'h3caa, 16'h3054,
// 16'h2307, 16'h14ff, 16'h0692, 16'hf7fa,
// 16'he994, 16'hdb99, 16'hce67, 16'hc227,
// 16'hb73a, 16'hadb2, 16'ha5eb, 16'h9fe1,
// 16'h9be0, 16'h99d1, 16'h99e6, 16'h9c20,
// 16'ha029, 16'ha63d, 16'hae2b, 16'hb7b4,
// 16'hc2c5, 16'hcf05, 16'hdc4b, 16'hea49,
// 16'hf8b5, 16'h074a, 16'h15b9, 16'h23b3,
// 16'h30fc, 16'h3d3c, 16'h484b, 16'h51d5,
// 16'h59c4, 16'h5fd6, 16'h6420, 16'h661c,
// 16'h662c, 16'h6423, 16'h601c, 16'h5a18,
// 16'h524b, 16'h48c9, 16'h3dd6, 16'h319a,
// 16'h2467, 16'h166c, 16'h0806, 16'hf96f,
// 16'heaff, 16'hdcfb, 16'hcfa9, 16'hc35a,
// 16'hb83a, 16'hae9c, 16'ha695, 16'ha06d,
// 16'h9c29, 16'h99f4, 16'h99c7, 16'h9bb6,
// 16'h9fa5, 16'ha58f, 16'had48, 16'hb6b3,
// 16'hc196, 16'hcdc1, 16'hdaed, 16'he8dc,
// 16'hf742, 16'h05d5, 16'h144a, 16'h2256,
// 16'h2fb0, 16'h3c13, 16'h473c, 16'h50f7,
// 16'h5909, 16'h5f56, 16'h63a7, 16'h6602,
// 16'h663e, 16'h6473, 16'h6096, 16'h5acc,
// 16'h5323, 16'h49d1, 16'h3efb, 16'h32e3,
// 16'h25c0, 16'h17da, 16'h097a, 16'hfae2,
// 16'hec70, 16'hde58, 16'hd0f6, 16'hc487,
// 16'hb947, 16'haf80, 16'ha74e, 16'ha0f5,
// 16'h9c7f, 16'h9a14, 16'h99b5, 16'h9b6b,
// 16'h9f2b, 16'ha4e1, 16'hac6e, 16'hb5b0,
// 16'hc070, 16'hcc7d, 16'hd992, 16'he771,
// 16'hf5cd, 16'h0461, 16'h12db, 16'h20f6,
// 16'h2e63, 16'h3ae3, 16'h462f, 16'h500f,
// 16'h5850, 16'h5ec8, 16'h6352, 16'h65db,
// 16'h6653, 16'h64b5, 16'h6114, 16'h5b72,
// 16'h53fd, 16'h4ad2, 16'h401f, 16'h3428,
// 16'h2717, 16'h1947, 16'h0aeb, 16'hfc5b,
// 16'heddc, 16'hdfbb, 16'hd242, 16'hc5b9,
// 16'hba58, 16'hb067, 16'ha80e, 16'ha17f,
// 16'h9cde, 16'h9a37, 16'h99a8, 16'h9b29,
// 16'h9eb2, 16'ha43a, 16'hab98, 16'hb4b1,
// 16'hbf4e, 16'hcb3a, 16'hd839, 16'he607,
// 16'hf45a, 16'h02ec, 16'h116b, 16'h1f93,
// 16'h2d17, 16'h39ad, 16'h4520, 16'h4f22,
// 16'h5792, 16'h5e37, 16'h62f5, 16'h65b3,
// 16'h665d, 16'h64f8, 16'h6186, 16'h5c19,
// 16'h54d1, 16'h4bcd, 16'h4143, 16'h3566,
// 16'h2871, 16'h1aaf, 16'h0c5e, 16'hfdd1,
// 16'hef4b, 16'he120, 16'hd391, 16'hc6ec,
// 16'hbb6e, 16'hb152, 16'ha8d1, 16'ha212,
// 16'h9d3a, 16'h9a68, 16'h999a, 16'h9aee,
// 16'h9e3e, 16'ha397, 16'haac9, 16'hb3b2,
// 16'hbe31, 16'hc9f9, 16'hd6e4, 16'he49e,
// 16'hf2e6, 16'h0178, 16'h0ffa, 16'h1e2f,
// 16'h2bc6, 16'h3878, 16'h4408, 16'h4e36,
// 16'h56cc, 16'h5da4, 16'h6292, 16'h6582,
// 16'h6668, 16'h6530, 16'h61f9, 16'h5cb7,
// 16'h55a1, 16'h4cc7, 16'h4260, 16'h36a4,
// 16'h29c7, 16'h1c17, 16'h0dd1, 16'hff45,
// 16'hf0bd, 16'he284, 16'hd4e4, 16'hc823,
// 16'hbc84, 16'hb244, 16'ha997, 16'ha2a8,
// 16'h9da2, 16'h9a95, 16'h999a, 16'h9ab2,
// 16'h9dd2, 16'ha2fa, 16'ha9f8, 16'hb2c1,
// 16'hbd0f, 16'hc8c1, 16'hd58d, 16'he337,
// 16'hf175, 16'h2001, 16'h0e8a, 16'h1cc9,
// 16'h2a73, 16'h3740, 16'h42ee, 16'h4d43,
// 16'h5605, 16'h5d07, 16'h622f, 16'h654a,
// 16'h666b, 16'h6566, 16'h6262, 16'h5d55,
// 16'h566b, 16'h4dbb, 16'h437c, 16'h37dd,
// 16'h2b1c, 16'h1d7c, 16'h0f44, 16'h20ba,
// 16'hf22f, 16'he3ea, 16'hd637, 16'hc95e,
// 16'hbda0, 16'hb337, 16'haa63, 16'ha344,
// 16'h9e0c, 16'h9acb, 16'h999e, 16'h9a79,
// 16'h9d71, 16'ha25b, 16'ha933, 16'hb1cc,
// 16'hbbf7, 16'hc788, 16'hd43a, 16'he1d2,
// 16'hf004, 16'hfe8a, 16'h0d19, 16'h1b61,
// 16'h291f, 16'h3604, 16'h41d1, 16'h4c4c,
// 16'h5538, 16'h5c6a, 16'h61c0, 16'h6513,
// 16'h6665, 16'h6599, 16'h62c7, 16'h5deb,
// 16'h5732, 16'h4eab, 16'h4495, 16'h3912,
// 16'h2c70, 16'h1ee0, 16'h10b5, 16'h022e,
// 16'hf3a3, 16'he551, 16'hd78f, 16'hca9a,
// 16'hbebd, 16'hb433, 16'hab2f, 16'ha3e7,
// 16'h9e7a, 16'h9b09, 16'h99a0, 16'h9a51,
// 16'h9d08, 16'ha1ca, 16'ha86f, 16'hb0db,
// 16'hbae3, 16'hc652, 16'hd2e8, 16'he06f,
// 16'hee93, 16'hfd16, 16'h0ba3, 16'h19fd,
// 16'h27c3, 16'h34c9, 16'h40b0, 16'h4b51,
// 16'h5466, 16'h5bc8, 16'h614c, 16'h64d8,
// 16'h665a, 16'h65c5, 16'h6326, 16'h5e7f,
// 16'h57f2, 16'h4f9a, 16'h45a6, 16'h3a4a,
// 16'h2dbc, 16'h2046, 16'h1223, 16'h03a5,
// 16'hf516, 16'he6b9, 16'hd8e7, 16'hcbdc,
// 16'hbfdd, 16'hb530, 16'hac03, 16'ha48d,
// 16'h9eed, 16'h9b4c, 16'h99aa, 16'h9a28,
// 16'h9cac, 16'ha139, 16'ha7b0, 16'haff0,
// 16'hb9d1, 16'hc520, 16'hd199, 16'hdf0d,
// 16'hed22, 16'hfba2, 16'h0a31, 16'h1890,
// 16'h266d, 16'h3384, 16'h3f91, 16'h4a4f,
// 16'h5391, 16'h5b20, 16'h60d4, 16'h6498,
// 16'h6647, 16'h65ef, 16'h637e, 16'h5f0f,
// 16'h58ad, 16'h5085, 16'h46b4, 16'h3b7d,
// 16'h2f08, 16'h21a8, 16'h1391, 16'h051c,
// 16'hf688, 16'he824, 16'hda43, 16'hcd1a,
// 16'hc107, 16'hb62d, 16'hacde, 16'ha535,
// 16'h9f69, 16'h9b8f, 16'h99be, 16'h9a03,
// 16'h9c54, 16'ha0ae, 16'ha6f5, 16'haf09,
// 16'hb8c5, 16'hc3eb, 16'hd053, 16'hdda8,
// 16'hebb6, 16'hfa2c, 16'h08bc, 16'h1726,
// 16'h2511, 16'h3241, 16'h3e68, 16'h494e,
// 16'h52b7, 16'h5a72, 16'h605b, 16'h644a,
// 16'h6637, 16'h660f, 16'h63d4, 16'h5f98,
// 16'h5965, 16'h5169, 16'h47c1, 16'h3cab,
// 16'h3053, 16'h2308, 16'h14ff, 16'h0691,
// 16'hf7fb, 16'he993, 16'hdb9b, 16'hce63,
// 16'hc22d, 16'hb733, 16'hadba, 16'ha5e4,
// 16'h9fe7, 16'h9bda, 16'h99d6, 16'h99e2,
// 16'h9c04, 16'ha025, 16'ha641, 16'hae26,
// 16'hb7ba, 16'hc2bf, 16'hcf09, 16'hdc49,
// 16'hea49, 16'hf8b6, 16'h074a, 16'h15b8,
// 16'h23b5, 16'h30f9, 16'h3d3f, 16'h4847,
// 16'h51da, 16'h59bf, 16'h5fdb, 16'h63fb,
// 16'h6620, 16'h6628, 16'h6428, 16'h6017,
// 16'h5a1c, 16'h5248, 16'h48ca, 16'h3dd6,
// 16'h319c, 16'h2463, 16'h1670, 16'h0802,
// 16'hf972, 16'heafe, 16'hdcfa, 16'hcfac,
// 16'hc356, 16'hb83e, 16'hae99, 16'ha697,
// 16'ha06d, 16'h9c28, 16'h99f3, 16'h99c9,
// 16'h9bb5, 16'h9fa6, 16'ha58e, 16'had47,
// 16'hb6b4, 16'hc196, 16'hcdc2, 16'hdaec,
// 16'he8dd, 16'hf740, 16'h05d7, 16'h1449,
// 16'h2257, 16'h2fb0, 16'h3c12, 16'h473c,
// 16'h50f8, 16'h5908, 16'h5f57, 16'h63a7,
// 16'h6620, 16'h6641, 16'h6471, 16'h6098,
// 16'h5ac9, 16'h5325, 16'h49cf, 16'h3efe,
// 16'h32e2, 16'h25be, 16'h17dd, 16'h0975,
// 16'hfae9, 16'hec6a, 16'hde5c, 16'hd0f4,
// 16'hc487, 16'hb948, 16'haf7f, 16'ha750,
// 16'ha0f3, 16'h9c81, 16'h9a12, 16'h99b5,
// 16'h9b6e, 16'h9f27, 16'ha4e5, 16'hac6b,
// 16'hb5b2, 16'hc06e, 16'hcc7e, 16'hd993,
// 16'he76e, 16'hf5d2, 16'h045b, 16'h12e0,
// 16'h20f2, 16'h2e66, 16'h3ae2, 16'h462e,
// 16'h5010, 16'h5850, 16'h5ec7, 16'h6353,
// 16'h65db, 16'h6651, 16'h64b9, 16'h6110,
// 16'h5b75, 16'h53fb, 16'h4ad2, 16'h4021,
// 16'h3425, 16'h271b, 16'h1943, 16'h0aed,
// 16'hfc5b, 16'hedda, 16'hdfbe, 16'hd240,
// 16'hc5ba, 16'hba57, 16'hb067, 16'ha80e,
// 16'ha180, 16'h9cdc, 16'h9a3a, 16'h99a5,
// 16'h9b29, 16'h9eb4, 16'ha438, 16'hab9a,
// 16'hb4b1, 16'hbf4b, 16'hcb3d, 16'hd838,
// 16'he607, 16'hf45b, 16'h02eb, 16'h116b,
// 16'h1f93, 16'h2d17, 16'h39ae, 16'h451e,
// 16'h4f23, 16'h5792, 16'h5e37, 16'h62f5,
// 16'h65b3, 16'h665c, 16'h64fa, 16'h6184,
// 16'h5c1b, 16'h54ce, 16'h4bd0, 16'h4141,
// 16'h3567, 16'h2871, 16'h1aaf, 16'h0c5e,
// 16'hfdd0, 16'hef4c, 16'he11f, 16'hd393,
// 16'hc6eb, 16'hbb6d, 16'hb153, 16'ha8d0,
// 16'ha212, 16'h9d3d, 16'h9a63, 16'h99a0,
// 16'h9ae7, 16'h9e44, 16'ha395, 16'haac7,
// 16'hb3b6, 16'hbe2d, 16'hc9fc, 16'hd6e3,
// 16'he49e, 16'hf2e6, 16'h0178, 16'h0ffa,
// 16'h1e2f, 16'h2bc7, 16'h3877, 16'h4409,
// 16'h4e34, 16'h56ce, 16'h5da3, 16'h6291,
// 16'h6585, 16'h6663, 16'h6535, 16'h61f4,
// 16'h5cbc, 16'h559c, 16'h4ccb, 16'h425d,
// 16'h36a6, 16'h29c5, 16'h1c19, 16'h0dce,
// 16'hff49, 16'hf0b9, 16'he288, 16'hd4e0,
// 16'hc825, 16'hbc84, 16'hb243, 16'ha999,
// 16'ha2a7, 16'h9da2, 16'h9a95, 16'h999a,
// 16'h9ab2, 16'h9dd3, 16'ha2f8, 16'ha9fb,
// 16'hb2bd, 16'hbd13, 16'hc8be, 16'hd58f,
// 16'he336, 16'hf175, 16'h2001, 16'h0e8a,
// 16'h1cc9, 16'h2a74, 16'h373d, 16'h42f2,
// 16'h4d40, 16'h5605, 16'h5d0b, 16'h6228,
// 16'h6552, 16'h6664, 16'h656b, 16'h6260,
// 16'h5d55, 16'h566b, 16'h4dbb, 16'h437c,
// 16'h37dd, 16'h2b1b, 16'h1d7f, 16'h0f40,
// 16'h20be, 16'hf22b, 16'he3ed, 16'hd636,
// 16'hc95f, 16'hbd9e, 16'hb33a, 16'haa60,
// 16'ha346, 16'h9e0b, 16'h9acc, 16'h999c,
// 16'h9a7c, 16'h9d6e, 16'ha25c, 16'ha934,
// 16'hb1ca, 16'hbbfa, 16'hc784, 16'hd43e,
// 16'he1cd, 16'hf008, 16'hfe89, 16'h0d18,
// 16'h1b63, 16'h291c, 16'h3606, 16'h41d0,
// 16'h4c4e, 16'h5535, 16'h5c6d, 16'h61bd,
// 16'h6516, 16'h6664, 16'h6599, 16'h62c6,
// 16'h5ded, 16'h5730, 16'h4eae, 16'h4491,
// 16'h3916, 16'h2c6c, 16'h1ee4, 16'h10b1,
// 16'h0233, 16'hf39f, 16'he552, 16'hd78f,
// 16'hca9a, 16'hbebd, 16'hb434, 16'hab2d,
// 16'ha3ea, 16'h9e77, 16'h9b0a, 16'h99a1,
// 16'h9a4f, 16'h9d0a, 16'ha1ca, 16'ha86d,
// 16'hb0dd, 16'hbae3, 16'hc650, 16'hd2ec,
// 16'he06b, 16'hee95, 16'hfd15, 16'h0ba5,
// 16'h19fb, 16'h27c4, 16'h34c8, 16'h40b0,
// 16'h4b53, 16'h5463, 16'h5bcb, 16'h6148,
// 16'h64dd, 16'h6654, 16'h65cb, 16'h6321,
// 16'h5e82, 16'h57f2, 16'h4f98, 16'h45a8,
// 16'h3a49, 16'h2dbc, 16'h2047, 16'h1222,
// 16'h03a5, 16'hf517, 16'he6b8, 16'hd8e9,
// 16'hcbd9, 16'hbfdf, 16'hb52f, 16'hac04,
// 16'ha48b, 16'h9ef1, 16'h9b46, 16'h99b0,
// 16'h9a24, 16'h9cad, 16'ha13b, 16'ha7ad,
// 16'haff2, 16'hb9d2, 16'hc51c, 16'hd19e,
// 16'hdf09, 16'hed25, 16'hfba0, 16'h0a32,
// 16'h1890, 16'h266c, 16'h3386, 16'h3f8e,
// 16'h4a50, 16'h5393, 16'h5b1e, 16'h60d5,
// 16'h6497, 16'h6647, 16'h65f0, 16'h637e,
// 16'h5f0e, 16'h58ae, 16'h5084, 16'h46b6,
// 16'h3b7a, 16'h2f0c, 16'h21a4, 16'h1394,
// 16'h051a, 16'hf689, 16'he825, 16'hda41,
// 16'hcd1d, 16'hc102, 16'hb633, 16'hacd9,
// 16'ha538, 16'h9f68, 16'h9b8d, 16'h99c2,
// 16'h99ff, 16'h9c57, 16'ha0ab, 16'ha6f8,
// 16'haf07, 16'hb8c7, 16'hc3ea, 16'hd052,
// 16'hdda9, 16'hebb6, 16'hfa2b, 16'h08bf,
// 16'h1722, 16'h2514, 16'h323f, 16'h3e69,
// 16'h494f, 16'h52b5, 16'h5a75, 16'h6056,
// 16'h6450, 16'h6633, 16'h6611, 16'h63d4,
// 16'h5f95, 16'h5969, 16'h5165, 16'h47c5,
// 16'h3ca8, 16'h3055, 16'h2306, 16'h1501,
// 16'h0690, 16'hf7fb, 16'he994, 16'hdb99,
// 16'hce66, 16'hc22a, 16'hb735, 16'hadb9,
// 16'ha5e4, 16'h9fe7, 16'h9bdb, 16'h99d5,
// 16'h99e3, 16'h9c02, 16'ha028, 16'ha63e,
// 16'hae29, 16'hb7b7, 16'hc2c2, 16'hcf05,
// 16'hdc4d, 16'hea46, 16'hf8b8, 16'h0749,
// 16'h15b8, 16'h23b5, 16'h30f9, 16'h3d3e,
// 16'h484a, 16'h51d7, 16'h59c1, 16'h5fd9,
// 16'h63fd, 16'h661e, 16'h662b, 16'h6424,
// 16'h601b, 16'h5a19, 16'h5249, 16'h48cc,
// 16'h3dd3, 16'h319f, 16'h2461, 16'h1671,
// 16'h0802, 16'hf971, 16'heb01, 16'hdcf6,
// 16'hcfaf, 16'hc354, 16'hb840, 16'hae97,
// 16'ha69a, 16'ha068, 16'h9c2d, 16'h99f0,
// 16'h99cc, 16'h9bb2, 16'h9fa8, 16'ha58c,
// 16'had4a, 16'hb6b2, 16'hc196, 16'hcdc3,
// 16'hdaeb, 16'he8dd, 16'hf742, 16'h05d4,
// 16'h144c, 16'h2254, 16'h2fb3, 16'h3c0f,
// 16'h473f, 16'h50f5, 16'h590b, 16'h5f53,
// 16'h63ab, 16'h65fd, 16'h6643, 16'h6470,
// 16'h6098, 16'h5aca, 16'h5324, 16'h49d0,
// 16'h3efd, 16'h32e2, 16'h25c0, 16'h17db,
// 16'h0977, 16'hfae6, 16'hec6d, 16'hde5a,
// 16'hd0f6, 16'hc485, 16'hb94a, 16'haf7c,
// 16'ha754, 16'ha0f0, 16'h9c82, 16'h9a12,
// 16'h99b5, 16'h9b6e, 16'h9f28, 16'ha4e3,
// 16'hac6c, 16'hb5b1, 16'hc071, 16'hcc7b,
// 16'hd994, 16'he76f, 16'hf5ce, 16'h0461,
// 16'h12da, 16'h20f7, 16'h2e63, 16'h3ae3,
// 16'h462e, 16'h500f, 16'h5851, 16'h5ec7,
// 16'h6353, 16'h65db, 16'h6651, 16'h64b8,
// 16'h6112, 16'h5b73, 16'h53fd, 16'h4ad0,
// 16'h4023, 16'h3422, 16'h271e, 16'h1941,
// 16'h0aef, 16'hfc58, 16'hedde, 16'hdfb9,
// 16'hd246, 16'hc5b4, 16'hba5b, 16'hb066,
// 16'ha80e, 16'ha181, 16'h9cdb, 16'h9a39,
// 16'h99a7, 16'h9b28, 16'h9eb4, 16'ha439,
// 16'hab98, 16'hb4b2, 16'hbf4c, 16'hcb3c,
// 16'hd839, 16'he605, 16'hf45d, 16'h02e9,
// 16'h116e, 16'h1f91, 16'h2d17, 16'h39ae,
// 16'h451f, 16'h4f22, 16'h5792, 16'h5e37,
// 16'h62f5, 16'h65b3, 16'h665d, 16'h64f8,
// 16'h6186, 16'h5c1a, 16'h54cf, 16'h4bcf,
// 16'h4142, 16'h3566, 16'h2871, 16'h1ab0,
// 16'h0c5d, 16'hfdd1, 16'hef4b, 16'he120,
// 16'hd391, 16'hc6ec, 16'hbb6e, 16'hb151,
// 16'ha8d2, 16'ha211, 16'h9d3c, 16'h9a66,
// 16'h999c, 16'h9aeb, 16'h9e40, 16'ha397,
// 16'haac8, 16'hb3b5, 16'hbe2e, 16'hc9fa,
// 16'hd6e4, 16'he49d, 16'hf2e9, 16'h0174,
// 16'h0ffe, 16'h1e2b, 16'h2bca, 16'h3874,
// 16'h440c, 16'h4e32, 16'h56d0, 16'h5da0,
// 16'h6295, 16'h6580, 16'h6669, 16'h6530,
// 16'h61f7, 16'h5cba, 16'h559e, 16'h4cc9,
// 16'h4260, 16'h36a2, 16'h29c9, 16'h1c15,
// 16'h0dd2, 16'hff46, 16'hf0bc, 16'he284,
// 16'hd4e3, 16'hc824, 16'hbc84, 16'hb244,
// 16'ha996, 16'ha2aa, 16'h9d9f, 16'h9a99,
// 16'h9996, 16'h9ab4, 16'h9dd3, 16'ha2f7,
// 16'ha9fc, 16'hb2be, 16'hbd10, 16'hc8c2,
// 16'hd58b, 16'he338, 16'hf176, 16'hffff,
// 16'h0e8c, 16'h1cc7, 16'h2a75, 16'h373d,
// 16'h42f2, 16'h4d40, 16'h5606, 16'h5d08,
// 16'h622c, 16'h654e, 16'h6668, 16'h6568,
// 16'h6261, 16'h5d56, 16'h5669, 16'h4dbe,
// 16'h4379, 16'h37df, 16'h2b1c, 16'h1d7b,
// 16'h0f45, 16'h20b9, 16'hf22f, 16'he3eb,
// 16'hd636, 16'hc95f, 16'hbd9e, 16'hb33a,
// 16'haa5f, 16'ha349, 16'h9e06, 16'h9ad1,
// 16'h9998, 16'h9a7f, 16'h9d6d, 16'ha25c,
// 16'ha935, 16'hb1c8, 16'hbbfb, 16'hc786,
// 16'hd43a, 16'he1d3, 16'hf001, 16'hfe8d,
// 16'h0d17, 16'h1b63, 16'h291d, 16'h3605,
// 16'h41d0, 16'h4c4d, 16'h5537, 16'h5c6b,
// 16'h61bf, 16'h6515, 16'h6663, 16'h659b,
// 16'h62c4, 16'h5dee, 16'h5731, 16'h4eaa,
// 16'h4497, 16'h3911, 16'h2c6f, 16'h1ee3,
// 16'h10b1, 16'h0232, 16'hf3a1, 16'he551,
// 16'hd790, 16'hca98, 16'hbec0, 16'hb42f,
// 16'hab34, 16'ha3e2, 16'h9e7e, 16'h9b06,
// 16'h99a2, 16'h9a4f, 16'h9d0b, 16'ha1c7,
// 16'ha872, 16'hb0d7, 16'hbae8, 16'hc64e,
// 16'hd2eb, 16'he06d, 16'hee93, 16'hfd16,
// 16'h0ba6, 16'h19f8, 16'h27c8, 16'h34c5,
// 16'h40b1, 16'h4b53, 16'h5463, 16'h5bcb,
// 16'h614a, 16'h64d9, 16'h6659, 16'h65c7,
// 16'h6324, 16'h5e81, 16'h57f1, 16'h4f9a,
// 16'h45a7, 16'h3a48, 16'h2dbe, 16'h2045,
// 16'h1223, 16'h03a6, 16'hf514, 16'he6bb,
// 16'hd8e6, 16'hcbdb, 16'hbfde, 16'hb530,
// 16'hac04, 16'ha48a, 16'h9ef1, 16'h9b46,
// 16'h99b0, 16'h9a24, 16'h9cae, 16'ha139,
// 16'ha7ae, 16'haff3, 16'hb9ce, 16'hc522,
// 16'hd198, 16'hdf0d, 16'hed24, 16'hfb9e,
// 16'h0a35, 16'h188d, 16'h266f, 16'h3384,
// 16'h3f8e, 16'h4a52, 16'h5390, 16'h5b21,
// 16'h60d3, 16'h6498, 16'h6646, 16'h65f1,
// 16'h637d, 16'h5f0f, 16'h58ad, 16'h5084,
// 16'h46b7, 16'h3b78, 16'h2f0e, 16'h21a2,
// 16'h1397, 16'h0518, 16'hf689, 16'he825,
// 16'hda42, 16'hcd1b, 16'hc107, 16'hb62c,
// 16'hacdf, 16'ha535, 16'h9f68, 16'h9b8f,
// 16'h99c0, 16'h9a20, 16'h9c57, 16'ha0ac,
// 16'ha6f6, 16'haf08, 16'hb8c6, 16'hc3eb,
// 16'hd053, 16'hdda7, 16'hebb8, 16'hfa29,
// 16'h08bf, 16'h1725, 16'h2511, 16'h3240,
// 16'h3e6a, 16'h494c, 16'h52b9, 16'h5a71,
// 16'h605a, 16'h644c, 16'h6637, 16'h660c,
// 16'h63d9, 16'h5f92, 16'h596a, 16'h5165,
// 16'h47c4, 16'h3ca9, 16'h3055, 16'h2306,
// 16'h1520, 16'h0691, 16'hf7fb, 16'he992,
// 16'hdb9d, 16'hce62, 16'hc22d, 16'hb733,
// 16'hadb9, 16'ha5e5, 16'h9fe7, 16'h9bda,
// 16'h99d5, 16'h99e4, 16'h9c01, 16'ha029,
// 16'ha63d, 16'hae29, 16'hb7b7, 16'hc2c2,
// 16'hcf07, 16'hdc4a, 16'hea49, 16'hf8b5,
// 16'h074b, 16'h15b7, 16'h23b6, 16'h30f8,
// 16'h3d40, 16'h4847, 16'h51da, 16'h59bf,
// 16'h5fda, 16'h63fd, 16'h661e, 16'h662a,
// 16'h6426, 16'h6018, 16'h5a1c, 16'h5247,
// 16'h48cc, 16'h3dd5, 16'h319b, 16'h2465,
// 16'h166e, 16'h0804, 16'hf972, 16'heafd,
// 16'hdcfa, 16'hcfad, 16'hc355, 16'hb840,
// 16'hae96, 16'ha69a, 16'ha06a, 16'h9c2b,
// 16'h99f1, 16'h99ca, 16'h9bb4, 16'h9fa6,
// 16'ha58f, 16'had47, 16'hb6b4, 16'hc195,
// 16'hcdc2, 16'hdaec, 16'he8de, 16'hf73f,
// 16'h05d9, 16'h1446, 16'h225a, 16'h2fad,
// 16'h3c14, 16'h473c, 16'h50f6, 16'h590c,
// 16'h5f51, 16'h63ad, 16'h65fc, 16'h6644,
// 16'h646e, 16'h609a, 16'h5ac9, 16'h5324,
// 16'h49d1, 16'h3efb, 16'h32e4, 16'h25bf,
// 16'h17da, 16'h0978, 16'hfae6, 16'hec6c,
// 16'hde5b, 16'hd0f5, 16'hc485, 16'hb94c,
// 16'haf7a, 16'ha754, 16'ha0f0, 16'h9c83,
// 16'h9a11, 16'h99b7, 16'h9b6b, 16'h9f2b,
// 16'ha4df, 16'hac72, 16'hb5ab, 16'hc075,
// 16'hcc79, 16'hd995, 16'he76f, 16'hf5cf,
// 16'h045f, 16'h12dc, 16'h20f6, 16'h2e63,
// 16'h3ae4, 16'h462d, 16'h5011, 16'h584f,
// 16'h5ec7, 16'h6354, 16'h65da, 16'h6653,
// 16'h64b6, 16'h6113, 16'h5b72, 16'h53ff,
// 16'h4ace, 16'h4024, 16'h3423, 16'h271b,
// 16'h1944, 16'h0aed, 16'hfc5a, 16'heddb,
// 16'hdfbe, 16'hd23f, 16'hc5bb, 16'hba56,
// 16'hb069, 16'ha80c, 16'ha182, 16'h9cda,
// 16'h9a3a, 16'h99a8, 16'h9b25, 16'h9eb7,
// 16'ha435, 16'hab9d, 16'hb4ae, 16'hbf4e,
// 16'hcb3b, 16'hd838, 16'he609, 16'hf458,
// 16'h02ed, 16'h116a, 16'h1f95, 16'h2d15,
// 16'h39af, 16'h451d, 16'h4f23, 16'h5794,
// 16'h5e35, 16'h62f6, 16'h65b1, 16'h665f,
// 16'h64f8, 16'h6185, 16'h5c1a, 16'h54cf,
// 16'h4bd0, 16'h4141, 16'h3567, 16'h2870,
// 16'h1ab0, 16'h0c5d, 16'hfdd2, 16'hef4a,
// 16'he120, 16'hd392, 16'hc6ea, 16'hbb70,
// 16'hb150, 16'ha8d3, 16'ha20f, 16'h9d3f,
// 16'h9a61, 16'h99a2, 16'h9ae7, 16'h9e43,
// 16'ha396, 16'haac5, 16'hb3b9, 16'hbe29,
// 16'hca01, 16'hd6de, 16'he4a0, 16'hf2e8,
// 16'h0174, 16'h0ffd, 16'h1e2e, 16'h2bc6,
// 16'h3879, 16'h4408, 16'h4e34, 16'h56cf,
// 16'h5da1, 16'h6295, 16'h6580, 16'h6667,
// 16'h6532, 16'h61f6, 16'h5cbb, 16'h559d,
// 16'h4cc9, 16'h425f, 16'h36a4, 16'h29c8,
// 16'h1c15, 16'h0dd2, 16'hff45, 16'hf0bd,
// 16'he285, 16'hd4e1, 16'hc826, 16'hbc82,
// 16'hb245, 16'ha997, 16'ha2a8, 16'h9da1,
// 16'h9a97, 16'h9998, 16'h9ab3, 16'h9dd3,
// 16'ha2f8, 16'ha9fb, 16'hb2be, 16'hbd11,
// 16'hc8c0, 16'hd58e, 16'he336, 16'hf177,
// 16'hffff, 16'h0e8a, 16'h1ccb, 16'h2a6f,
// 16'h3745, 16'h42ea, 16'h4d46, 16'h5602,
// 16'h5d0a, 16'h622b, 16'h6550, 16'h6665,
// 16'h656b, 16'h625f, 16'h5d56, 16'h566a,
// 16'h4dbd, 16'h4379, 16'h37e0, 16'h2b1a,
// 16'h1d7d, 16'h0f43, 16'h20bb, 16'hf22e,
// 16'he3eb, 16'hd637, 16'hc95e, 16'hbd9e,
// 16'hb33b, 16'haa5f, 16'ha347, 16'h9e0a,
// 16'h9acd, 16'h999b, 16'h9a7d, 16'h9d6d,
// 16'ha25e, 16'ha932, 16'hb1cc, 16'hbbf6,
// 16'hc789, 16'hd43a, 16'he1d1, 16'hf006,
// 16'hfe87, 16'h0d1b, 16'h1b60, 16'h2920,
// 16'h3603, 16'h41d2, 16'h4c4c, 16'h5536,
// 16'h5c6d, 16'h61bd, 16'h6517, 16'h6662,
// 16'h659a, 16'h62c6, 16'h5dec, 16'h5732,
// 16'h4eac, 16'h4492, 16'h3917, 16'h2c6a,
// 16'h1ee5, 16'h10b1, 16'h0233, 16'hf39f,
// 16'he553, 16'hd78d, 16'hca9b, 16'hbebe,
// 16'hb432, 16'hab2f, 16'ha3e8, 16'h9e78,
// 16'h9b0a, 16'h99a2, 16'h9a4c, 16'h9d0e,
// 16'ha1c5, 16'ha871, 16'hb0dc, 16'hbae2,
// 16'hc651, 16'hd2eb, 16'he06c, 16'hee94,
// 16'hfd16, 16'h0ba5, 16'h19f9, 16'h27c9,
// 16'h34c2, 16'h40b5, 16'h4b4f, 16'h5467,
// 16'h5bc7, 16'h614e, 16'h64d5, 16'h665d,
// 16'h65c2, 16'h6329, 16'h5e7c, 16'h57f5,
// 16'h4f98, 16'h45a6, 16'h3a4b, 16'h2dbb,
// 16'h2047, 16'h1221, 16'h03a8, 16'hf512,
// 16'he6be, 16'hd8e3, 16'hcbdd, 16'hbfdd,
// 16'hb531, 16'hac02, 16'ha48c, 16'h9ef0,
// 16'h9b47, 16'h99af, 16'h9a26, 16'h9caa,
// 16'ha13d, 16'ha7ac, 16'haff3, 16'hb9d0,
// 16'hc51e, 16'hd19c, 16'hdf0b, 16'hed24,
// 16'hfba0, 16'h0a31, 16'h1891, 16'h266c,
// 16'h3385, 16'h3f90, 16'h4a4e, 16'h5394,
// 16'h5b1d, 16'h60d7, 16'h6494, 16'h664a,
// 16'h65ee, 16'h637f, 16'h5f0e, 16'h58ae,
// 16'h5083, 16'h46b6, 16'h3b7c, 16'h2f08,
// 16'h21aa, 16'h138f, 16'h051e, 16'hf685,
// 16'he828, 16'hda3f, 16'hcd1f, 16'hc103,
// 16'hb630, 16'hacdb, 16'ha538, 16'h9f65,
// 16'h9b93, 16'h99bc, 16'h9a03, 16'h9c54,
// 16'ha0ae, 16'ha6f5, 16'haf0a, 16'hb8c4,
// 16'hc3eb, 16'hd054, 16'hdda7, 16'hebb7,
// 16'hfa2a, 16'h08bf, 16'h1724, 16'h2513,
// 16'h323f, 16'h3e69, 16'h494e, 16'h52b6,
// 16'h5a74, 16'h6059, 16'h644c, 16'h6637,
// 16'h660d, 16'h63d6, 16'h5f96, 16'h5967,
// 16'h5168, 16'h47c2, 16'h3ca9, 16'h3055,
// 16'h2307, 16'h14ff, 16'h0692, 16'hf7f9,
// 16'he995, 16'hdb9a, 16'hce64, 16'hc22a,
// 16'hb738, 16'hadb4, 16'ha5e9, 16'h9fe4,
// 16'h9bda, 16'h99d8, 16'h99e0, 16'h9c05,
// 16'ha025, 16'ha641, 16'hae24, 16'hb7bd,
// 16'hc2bd, 16'hcf0b, 16'hdc47, 16'hea4b,
// 16'hf8b4, 16'h074b, 16'h15b8, 16'h23b5,
// 16'h30f8, 16'h3d41, 16'h4845, 16'h51db,
// 16'h59bf, 16'h5fda, 16'h63fc, 16'h661f,
// 16'h6629, 16'h6426, 16'h601a, 16'h5a1a,
// 16'h5248, 16'h48cb, 16'h3dd5, 16'h319c,
// 16'h2465, 16'h166e, 16'h0802, 16'hf974,
// 16'heafb, 16'hdcfd, 16'hcfaa, 16'hc357,
// 16'hb83e, 16'hae97, 16'ha69b, 16'ha067,
// 16'h9c2f, 16'h99ed, 16'h99ce, 16'h9bb1,
// 16'h9fa8, 16'ha58e, 16'had46, 16'hb6b6,
// 16'hc194, 16'hcdc3, 16'hdaec, 16'he8dc,
// 16'hf742, 16'h05d5, 16'h144c, 16'h2253,
// 16'h2fb3, 16'h3c10, 16'h473e, 16'h50f6,
// 16'h590c, 16'h5f50, 16'h63ae, 16'h65fb,
// 16'h6644, 16'h6470, 16'h6097, 16'h5acc,
// 16'h5322, 16'h49d2, 16'h3efb, 16'h32e2,
// 16'h25c1, 16'h17da, 16'h0977, 16'hfae7,
// 16'hec6c, 16'hde59, 16'hd0f8, 16'hc482,
// 16'hb94d, 16'haf7b, 16'ha753, 16'ha0f1,
// 16'h9c82, 16'h9a12, 16'h99b6, 16'h9b6c,
// 16'h9f29, 16'ha4e2, 16'hac6f, 16'hb5af,
// 16'hc071, 16'hcc7c, 16'hd990, 16'he775,
// 16'hf5c9, 16'h0466, 16'h12d6, 16'h20fa,
// 16'h2e5f, 16'h3ae7, 16'h462c, 16'h5011,
// 16'h5850, 16'h5ec6, 16'h6354, 16'h65da,
// 16'h6654, 16'h64b4, 16'h6115, 16'h5b71,
// 16'h53fe, 16'h4ad1, 16'h4020, 16'h3427,
// 16'h2718, 16'h1946, 16'h0aeb, 16'hfc5c,
// 16'heddb, 16'hdfbb, 16'hd243, 16'hc5b7,
// 16'hba5a, 16'hb065, 16'ha810, 16'ha17e,
// 16'h9cde, 16'h9a36, 16'h99aa, 16'h9b26,
// 16'h9eb4, 16'ha43b, 16'hab95, 16'hb4b5,
// 16'hbf49, 16'hcb3e, 16'hd838, 16'he606,
// 16'hf45d, 16'h02e8, 16'h116e, 16'h1f93,
// 16'h2d14, 16'h39b2, 16'h451a, 16'h4f27,
// 16'h578f, 16'h5e39, 16'h62f4, 16'h65b2,
// 16'h665e, 16'h64f9, 16'h6184, 16'h5c1b,
// 16'h54cf, 16'h4bcf, 16'h4142, 16'h3565,
// 16'h2872, 16'h1aaf, 16'h0c5e, 16'hfdd1,
// 16'hef4b, 16'he11f, 16'hd392, 16'hc6ec,
// 16'hbb6c, 16'hb155, 16'ha8ce, 16'ha214,
// 16'h9d3b, 16'h9a64, 16'h99a0, 16'h9ae7,
// 16'h9e44, 16'ha394, 16'haac9, 16'hb3b5,
// 16'hbe2c, 16'hc9ff, 16'hd6de, 16'he4a3,
// 16'hf2e4, 16'h0178, 16'h0ff9, 16'h1e32,
// 16'h2bc2, 16'h387d, 16'h4404, 16'h4e38,
// 16'h56cb, 16'h5da4, 16'h6292, 16'h6583,
// 16'h6666, 16'h6532, 16'h61f6, 16'h5cb9,
// 16'h55a1, 16'h4cc5, 16'h4263, 16'h36a1,
// 16'h29c8, 16'h1c17, 16'h0dd0, 16'hff46,
// 16'hf0bd, 16'he284, 16'hd4e3, 16'hc824,
// 16'hbc84, 16'hb243, 16'ha998, 16'ha2a9,
// 16'h9da0, 16'h9a97, 16'h9999, 16'h9ab0,
// 16'h9dd8, 16'ha2f4, 16'ha9fc, 16'hb2be,
// 16'hbd11, 16'hc8c1, 16'hd58d, 16'he336,
// 16'hf176, 16'h2001, 16'h0e8a, 16'h1cc9,
// 16'h2a73, 16'h373f, 16'h42f0, 16'h4d42,
// 16'h5605, 16'h5d08, 16'h622d, 16'h654c,
// 16'h666b, 16'h6566, 16'h6261, 16'h5d57,
// 16'h5667, 16'h4dc0, 16'h4379, 16'h37de,
// 16'h2b1c, 16'h1d7b, 16'h0f45, 16'h20b9,
// 16'hf230, 16'he3e9, 16'hd639, 16'hc95b,
// 16'hbda2, 16'hb337, 16'haa62, 16'ha346,
// 16'h9e09, 16'h9ace, 16'h999a, 16'h9a7e,
// 16'h9d6d, 16'ha25e, 16'ha931, 16'hb1cc,
// 16'hbbf8, 16'hc787, 16'hd43c, 16'he1ce,
// 16'hf008, 16'hfe87, 16'h0d1b, 16'h1b61,
// 16'h291d, 16'h3605, 16'h41d1, 16'h4c4c,
// 16'h5538, 16'h5c6b, 16'h61bd, 16'h6517,
// 16'h6661, 16'h659d, 16'h62c3, 16'h5def,
// 16'h572f, 16'h4ead, 16'h4493, 16'h3915,
// 16'h2c6c, 16'h1ee5, 16'h10b0, 16'h0234,
// 16'hf39c, 16'he558, 16'hd788, 16'hcaa0,
// 16'hbeb9, 16'hb435, 16'hab2e, 16'ha3e9,
// 16'h9e77, 16'h9b0b, 16'h999f, 16'h9a51,
// 16'h9d09, 16'ha1ca, 16'ha86d, 16'hb0de,
// 16'hbae1, 16'hc652, 16'hd2ea, 16'he06c,
// 16'hee96, 16'hfd13, 16'h0ba7, 16'h19f9,
// 16'h27c6, 16'h34c7, 16'h40b0, 16'h4b52,
// 16'h5466, 16'h5bc7, 16'h614d, 16'h64d8,
// 16'h6658, 16'h65c8, 16'h6323, 16'h5e82,
// 16'h57f0, 16'h4f9c, 16'h45a4, 16'h3a4b,
// 16'h2dbc, 16'h2045, 16'h1225, 16'h03a4,
// 16'hf516, 16'he6b9, 16'hd8e8, 16'hcbd9,
// 16'hbfe0, 16'hb52f, 16'hac03, 16'ha48d,
// 16'h9eed, 16'h9b4b, 16'h99ac, 16'h9a26,
// 16'h9cae, 16'ha137, 16'ha7b1, 16'haff1,
// 16'hb9d0, 16'hc51f, 16'hd19b, 16'hdf0b,
// 16'hed24, 16'hfba0, 16'h0a32, 16'h1890,
// 16'h266d, 16'h3384, 16'h3f8f, 16'h4a51,
// 16'h5391, 16'h5b20, 16'h60d5, 16'h6495,
// 16'h664a, 16'h65ed, 16'h6380, 16'h5f0d,
// 16'h58b0, 16'h5081, 16'h46b8, 16'h3b79,
// 16'h2f0c, 16'h21a5, 16'h1394, 16'h0519,
// 16'hf68a, 16'he823, 16'hda44, 16'hcd1a,
// 16'hc106, 16'hb62f, 16'hacda, 16'ha53a,
// 16'h9f64, 16'h9b93, 16'h99bc, 16'h9a03,
// 16'h9c55, 16'ha0ad, 16'ha6f6, 16'haf09,
// 16'hb8c4, 16'hc3ec, 16'hd054, 16'hdda5,
// 16'hebbb, 16'hfa26, 16'h08c1, 16'h1723,
// 16'h2513, 16'h3240, 16'h3e68, 16'h494f,
// 16'h52b5, 16'h5a75, 16'h6058, 16'h644c,
// 16'h6637, 16'h660e, 16'h63d5, 16'h5f96,
// 16'h5968, 16'h5166, 16'h47c4, 16'h3ca8,
// 16'h3056, 16'h2305, 16'h1501, 16'h0691,
// 16'hf7fa, 16'he994, 16'hdb9a, 16'hce65,
// 16'hc22a, 16'hb737, 16'hadb6, 16'ha5e6,
// 16'h9fe6, 16'h9bdb, 16'h99d6, 16'h99e1,
// 16'h9c04, 16'ha026, 16'ha640, 16'hae27,
// 16'hb7b9, 16'hc2bf, 16'hcf0a, 16'hdc48,
// 16'hea4a, 16'hf8b6, 16'h0748, 16'h15bb,
// 16'h23b2, 16'h30fb, 16'h3d3f, 16'h4846,
// 16'h51db, 16'h59be, 16'h5fdc, 16'h63fb,
// 16'h6620, 16'h6628, 16'h6427, 16'h6019,
// 16'h5a1a, 16'h5249, 16'h48cb, 16'h3dd4,
// 16'h319e, 16'h2462, 16'h1670, 16'h0802,
// 16'hf973, 16'heafc, 16'hdcfd, 16'hcfa8,
// 16'hc35a, 16'hb83b, 16'hae9a, 16'ha698,
// 16'ha06a, 16'h9c2c, 16'h99f0, 16'h99cb,
// 16'h9bb3, 16'h9fa7, 16'ha58e, 16'had48,
// 16'hb6b3, 16'hc197, 16'hcdbe, 16'hdaf2,
// 16'he8d7, 16'hf746, 16'h05d2, 16'h144c,
// 16'h2256, 16'h2fae, 16'h3c15, 16'h473b,
// 16'h50f7, 16'h590c, 16'h5f50, 16'h63ad,
// 16'h65fd, 16'h6643, 16'h646f, 16'h609a,
// 16'h5ac8, 16'h5325, 16'h49cf, 16'h3efe,
// 16'h32e0, 16'h25c3, 16'h17d8, 16'h0978,
// 16'hfae7, 16'hec6b, 16'hde5b, 16'hd0f6,
// 16'hc484, 16'hb94b, 16'haf7d, 16'ha750,
// 16'ha0f5, 16'h9c7d, 16'h9a16, 16'h99b4,
// 16'h9b6c, 16'h9f2b, 16'ha4df, 16'hac71,
// 16'hb5ae, 16'hc071, 16'hcc7c, 16'hd993,
// 16'he770, 16'hf5ce, 16'h0460, 16'h12dc,
// 16'h20f5, 16'h2e65, 16'h3ae1, 16'h4630,
// 16'h500f, 16'h584f, 16'h5eca, 16'h6350,
// 16'h65dd, 16'h6651, 16'h64b7, 16'h6112,
// 16'h5b73, 16'h53fe, 16'h4acf, 16'h4023,
// 16'h3423, 16'h271c, 16'h1944, 16'h0aec,
// 16'hfc5a, 16'heddd, 16'hdfbb, 16'hd243,
// 16'hc5b7, 16'hba59, 16'hb067, 16'ha80e,
// 16'ha17f, 16'h9cdd, 16'h9a37, 16'h99aa,
// 16'h9b25, 16'h9eb6, 16'ha436, 16'hab9c,
// 16'hb4ae, 16'hbf50, 16'hcb38, 16'hd83b,
// 16'he606, 16'hf45b, 16'h02eb, 16'h116c,
// 16'h1f93, 16'h2d15, 16'h39b0, 16'h451d,
// 16'h4f24, 16'h5792, 16'h5e35, 16'h62f8,
// 16'h65af, 16'h6660, 16'h64f7, 16'h6186,
// 16'h5c19, 16'h54d1, 16'h4bcd, 16'h4143,
// 16'h3566, 16'h2870, 16'h1ab1, 16'h0c5c,
// 16'hfdd2, 16'hef4b, 16'he120, 16'hd391,
// 16'hc6ec, 16'hbb6c, 16'hb155, 16'ha8cf,
// 16'ha213, 16'h9d3a, 16'h9a67, 16'h999c,
// 16'h9aeb, 16'h9e41, 16'ha395, 16'haaca,
// 16'hb3b2, 16'hbe30, 16'hc9fb, 16'hd6e3,
// 16'he49d, 16'hf2e9, 16'h0173, 16'h0fff,
// 16'h1e2d, 16'h2bc6, 16'h3878, 16'h440a,
// 16'h4e31, 16'h56d2, 16'h5d9f, 16'h6295,
// 16'h6583, 16'h6663, 16'h6536, 16'h61f2,
// 16'h5cbe, 16'h559d, 16'h4cc8, 16'h4260,
// 16'h36a3, 16'h29c8, 16'h1c16, 16'h0dd2,
// 16'hff43, 16'hf0c0, 16'he281, 16'hd4e6,
// 16'hc821, 16'hbc86, 16'hb243, 16'ha997,
// 16'ha2a9, 16'h9da0, 16'h9a98, 16'h9997,
// 16'h9ab4, 16'h9dd2, 16'ha2f9, 16'ha9f9,
// 16'hb2c0, 16'hbd0f, 16'hc8c3, 16'hd58a,
// 16'he33a, 16'hf172, 16'h2004, 16'h0e86,
// 16'h1cce, 16'h2a6e, 16'h3743, 16'h42ee,
// 16'h4d41, 16'h5607, 16'h5d07, 16'h622c,
// 16'h654f, 16'h6667, 16'h6569, 16'h6260,
// 16'h5d56, 16'h566a, 16'h4dbc, 16'h437c,
// 16'h37dd, 16'h2b1b, 16'h1d7e, 16'h0f41,
// 16'h20bc, 16'hf22f, 16'he3e9, 16'hd638,
// 16'hc95e, 16'hbd9d, 16'hb33c, 16'haa5e,
// 16'ha348, 16'h9e09, 16'h9ace, 16'h999a,
// 16'h9a7d, 16'h9d6e, 16'ha25c, 16'ha934,
// 16'hb1cb, 16'hbbf7, 16'hc788, 16'hd43a,
// 16'he1d1, 16'hf005, 16'hfe8a, 16'h0d18,
// 16'h1b63, 16'h291d, 16'h3605, 16'h41d0,
// 16'h4c4f, 16'h5532, 16'h5c72, 16'h61b8,
// 16'h651b, 16'h665f, 16'h659c, 16'h62c5,
// 16'h5dee, 16'h572f, 16'h4eaf, 16'h448f,
// 16'h3919, 16'h2c6a, 16'h1ee5, 16'h10b1,
// 16'h0231, 16'hf3a1, 16'he553, 16'hd78c,
// 16'hca9e, 16'hbeb9, 16'hb436, 16'hab2e,
// 16'ha3e7, 16'h9e7b, 16'h9b07, 16'h99a2,
// 16'h9a50, 16'h9d08, 16'ha1cb, 16'ha86e,
// 16'hb0db, 16'hbae5, 16'hc64e, 16'hd2ed,
// 16'he06b, 16'hee96, 16'hfd12, 16'h0ba8,
// 16'h19f8, 16'h27c8, 16'h34c5, 16'h40b1,
// 16'h4b52, 16'h5464, 16'h5bcb, 16'h6149,
// 16'h64db, 16'h6657, 16'h65c7, 16'h6325,
// 16'h5e7f, 16'h57f4, 16'h4f98, 16'h45a8,
// 16'h3a47, 16'h2dbf, 16'h2043, 16'h1226,
// 16'h03a4, 16'hf516, 16'he6b9, 16'hd8e7,
// 16'hcbda, 16'hbfe1, 16'hb52d, 16'hac05,
// 16'ha48a, 16'h9ef0, 16'h9b49, 16'h99ae,
// 16'h9a24, 16'h9cae, 16'ha139, 16'ha7af,
// 16'haff2, 16'hb9cf, 16'hc520, 16'hd19a,
// 16'hdf0d, 16'hed21, 16'hfba3, 16'h0a2f,
// 16'h1893, 16'h266a, 16'h3387, 16'h3f8c,
// 16'h4a54, 16'h538f, 16'h5b21, 16'h60d4,
// 16'h6495, 16'h664b, 16'h65ec, 16'h6382,
// 16'h5f0a, 16'h58b1, 16'h5082, 16'h46b6,
// 16'h3b7c, 16'h2f08, 16'h21a8, 16'h1391,
// 16'h051e, 16'hf684, 16'he829, 16'hda3e,
// 16'hcd1f, 16'hc102, 16'hb633, 16'hacd7,
// 16'ha53c, 16'h9f63, 16'h9b92, 16'h99be,
// 16'h9a01, 16'h9c57, 16'ha0aa, 16'ha6f9,
// 16'haf07, 16'hb8c5, 16'hc3ed, 16'hd04f,
// 16'hddac, 16'hebb3, 16'hfa2e, 16'h08bc,
// 16'h1726, 16'h2510, 16'h3242, 16'h3e67,
// 16'h4950, 16'h52b5, 16'h5a75, 16'h6057,
// 16'h644e, 16'h6634, 16'h6610, 16'h63d5,
// 16'h5f95, 16'h5969, 16'h5165, 16'h47c5,
// 16'h3ca8, 16'h3054, 16'h2308, 16'h1520,
// 16'h068f, 16'hf7fe, 16'he98f, 16'hdb9e,
// 16'hce63, 16'hc22b, 16'hb736, 16'hadb6,
// 16'ha5e6, 16'h9fe7, 16'h9bda, 16'h99d7,
// 16'h99e1, 16'h9c03, 16'ha027, 16'ha63f,
// 16'hae29, 16'hb7b6, 16'hc2c3, 16'hcf06,
// 16'hdc4a, 16'hea4b, 16'hf8b2, 16'h074e,
// 16'h15b4, 16'h23b9, 16'h30f6, 16'h3d41,
// 16'h4846, 16'h51da, 16'h59c0, 16'h5fda,
// 16'h63fc, 16'h661f, 16'h6629, 16'h6426,
// 16'h601a, 16'h5a19, 16'h524a, 16'h48ca,
// 16'h3dd5, 16'h319c, 16'h2465, 16'h166d,
// 16'h0806, 16'hf96e, 16'heb01, 16'hdcf9,
// 16'hcfab, 16'hc359, 16'hb83b, 16'hae9a,
// 16'ha698, 16'ha06a, 16'h9c2d, 16'h99ef,
// 16'h99cc, 16'h9bb1, 16'h9faa, 16'ha58b,
// 16'had4b, 16'hb6b0, 16'hc198, 16'hcdc0,
// 16'hdaee, 16'he8dc, 16'hf741, 16'h05d6,
// 16'h1449, 16'h2258, 16'h2fae, 16'h3c14,
// 16'h473b, 16'h50f8, 16'h5909, 16'h5f54,
// 16'h63ab, 16'h65fd, 16'h6643, 16'h646f,
// 16'h6099, 16'h5aca, 16'h5324, 16'h49d0,
// 16'h3efd, 16'h32e1, 16'h25c1, 16'h17db,
// 16'h0976, 16'hfae7, 16'hec6c, 16'hde5a,
// 16'hd0f6, 16'hc486, 16'hb948, 16'haf80,
// 16'ha74e, 16'ha0f4, 16'h9c81, 16'h9a12,
// 16'h99b6, 16'h9b6d, 16'h9f27, 16'ha4e5,
// 16'hac6b, 16'hb5b2, 16'hc06f, 16'hcc7e,
// 16'hd990, 16'he773, 16'hf5cd, 16'h045f,
// 16'h12de, 16'h20f3, 16'h2e65, 16'h3ae3,
// 16'h462d, 16'h5011, 16'h5850, 16'h5ec6,
// 16'h6355, 16'h65d8, 16'h6654, 16'h64b7,
// 16'h6110, 16'h5b76, 16'h53fa, 16'h4ad3,
// 16'h4020, 16'h3425, 16'h271b, 16'h1944,
// 16'h0aec, 16'hfc5b, 16'heddb, 16'hdfbd,
// 16'hd242, 16'hc5b7, 16'hba5a, 16'hb065,
// 16'ha80f, 16'ha180, 16'h9cdb, 16'h9a3b,
// 16'h99a4, 16'h9b2b, 16'h9eb0, 16'ha43d,
// 16'hab95, 16'hb4b4, 16'hbf4b, 16'hcb3b,
// 16'hd83b, 16'he604, 16'hf45d, 16'h02e9,
// 16'h116e, 16'h1f91, 16'h2d18, 16'h39ad,
// 16'h451f, 16'h4f22, 16'h5794, 16'h5e35,
// 16'h62f7, 16'h65b1, 16'h665d, 16'h64fa,
// 16'h6184, 16'h5c1b, 16'h54cf, 16'h4bce,
// 16'h4143, 16'h3565, 16'h2873, 16'h1aad,
// 16'h0c60, 16'hfdcf, 16'hef4c, 16'he120,
// 16'hd391, 16'hc6ec, 16'hbb6e, 16'hb151,
// 16'ha8d2, 16'ha211, 16'h9d3c, 16'h9a66,
// 16'h999b, 16'h9aee, 16'h9e3c, 16'ha39c,
// 16'haac2, 16'hb3b9, 16'hbe2c, 16'hc9fd,
// 16'hd6e1, 16'he49f, 16'hf2e7, 16'h0176,
// 16'h0ffb, 16'h1e30, 16'h2bc4, 16'h387a,
// 16'h4408, 16'h4e33, 16'h56d0, 16'h5da1,
// 16'h6293, 16'h6584, 16'h6663, 16'h6535,
// 16'h61f4, 16'h5cbb, 16'h55a0, 16'h4cc5,
// 16'h4263, 16'h36a1, 16'h29c9, 16'h1c16,
// 16'h0dd2, 16'hff44, 16'hf0bf, 16'he281,
// 16'hd4e6, 16'hc822, 16'hbc85, 16'hb244,
// 16'ha995, 16'ha2ab, 16'h9d9f, 16'h9a98,
// 16'h9998, 16'h9ab2, 16'h9dd4, 16'ha2f7,
// 16'ha9fc, 16'hb2be, 16'hbd10, 16'hc8c1,
// 16'hd58c, 16'he338, 16'hf176, 16'h2020,
// 16'h0e89, 16'h1ccb, 16'h2a70, 16'h3742,
// 16'h42ef, 16'h4d41, 16'h5605, 16'h5d0a,
// 16'h6229, 16'h6552, 16'h6664, 16'h656b,
// 16'h625f, 16'h5d56, 16'h566b, 16'h4dbb,
// 16'h437c, 16'h37dd, 16'h2b1c, 16'h1d7c,
// 16'h0f44, 16'h20b9, 16'hf231, 16'he3e8,
// 16'hd639, 16'hc95d, 16'hbda0, 16'hb337,
// 16'haa64, 16'ha343, 16'h9e0c, 16'h9acd,
// 16'h9999, 16'h9a80, 16'h9d6b, 16'ha25f,
// 16'ha931, 16'hb1cc, 16'hbbf8, 16'hc787,
// 16'hd43b, 16'he1d0, 16'hf006, 16'hfe89,
// 16'h0d1a, 16'h1b5f, 16'h2922, 16'h35ff,
// 16'h41d7, 16'h4c47, 16'h553b, 16'h5c69,
// 16'h61be, 16'h6517, 16'h6662, 16'h659b,
// 16'h62c5, 16'h5dec, 16'h5733, 16'h4eaa,
// 16'h4496, 16'h3911, 16'h2c71, 16'h1edf,
// 16'h10b6, 16'h022e, 16'hf3a3, 16'he550,
// 16'hd790, 16'hca99, 16'hbebe, 16'hb431,
// 16'hab31, 16'ha3e6, 16'h9e7b, 16'h9b07,
// 16'h99a3, 16'h9a4d, 16'h9d0c, 16'ha1c8,
// 16'ha86f, 16'hb0dd, 16'hbae0, 16'hc655,
// 16'hd2e6, 16'he071, 16'hee91, 16'hfd16,
// 16'h0ba5, 16'h19fa, 16'h27c6, 16'h34c7,
// 16'h40b0, 16'h4b52, 16'h5465, 16'h5bc9,
// 16'h614b, 16'h64d9, 16'h6658, 16'h65c8,
// 16'h6323, 16'h5e82, 16'h57ef, 16'h4f9d,
// 16'h45a3, 16'h3a4d, 16'h2db9, 16'h2049,
// 16'h1220, 16'h03a8, 16'hf514, 16'he6ba,
// 16'hd8e9, 16'hcbd6, 16'hbfe3, 16'hb52d,
// 16'hac04, 16'ha48c, 16'h9eee, 16'h9b4a,
// 16'h99ad, 16'h9a25, 16'h9cae, 16'ha137,
// 16'ha7b3, 16'hafed, 16'hb9d4, 16'hc51c,
// 16'hd19c, 16'hdf0d, 16'hed20, 16'hfba5,
// 16'h0a2d, 16'h1894, 16'h266a, 16'h3386,
// 16'h3f8d, 16'h4a55, 16'h538c, 16'h5b24,
// 16'h60d2, 16'h6495, 16'h664d, 16'h65ea,
// 16'h6382, 16'h5f0c, 16'h58af, 16'h5083,
// 16'h46b7, 16'h3b79, 16'h2f0c, 16'h21a6,
// 16'h1392, 16'h051c, 16'hf686, 16'he827,
// 16'hda40, 16'hcd1e, 16'hc103, 16'hb630,
// 16'hacdb, 16'ha537, 16'h9f68, 16'h9b8f,
// 16'h99bf, 16'h9a20, 16'h9c58, 16'ha0aa,
// 16'ha6f8, 16'haf08, 16'hb8c4, 16'hc3ee,
// 16'hd04f, 16'hddaa, 16'hebb6, 16'hfa2c,
// 16'h08bc, 16'h1726, 16'h2511, 16'h3241,
// 16'h3e68, 16'h494f, 16'h52b6, 16'h5a74,
// 16'h6057, 16'h644f, 16'h6633, 16'h6612,
// 16'h63d2, 16'h5f98, 16'h5965, 16'h516a,
// 16'h47c0, 16'h3cac, 16'h3052, 16'h2308,
// 16'h1520, 16'h068f, 16'hf7fe, 16'he98f,
// 16'hdb9f, 16'hce61, 16'hc22d, 16'hb734,
// 16'hadb7, 16'ha5e7, 16'h9fe5, 16'h9bdb,
// 16'h99d6, 16'h99e2, 16'h9c03, 16'ha027,
// 16'ha63f, 16'hae27, 16'hb7ba, 16'hc2bf,
// 16'hcf08, 16'hdc4b, 16'hea48, 16'hf8b7,
// 16'h0748, 16'h15b9, 16'h23b4, 16'h30fc,
// 16'h3d3c, 16'h4849, 16'h51d8, 16'h59c1,
// 16'h5fd9, 16'h63fe, 16'h661d, 16'h662a,
// 16'h6426, 16'h6019, 16'h5a1b, 16'h5248,
// 16'h48cc, 16'h3dd3, 16'h319e, 16'h2463,
// 16'h166e, 16'h0805, 16'hf970, 16'heaff,
// 16'hdcfa, 16'hcfab, 16'hc357, 16'hb83d,
// 16'hae9a, 16'ha696, 16'ha06e, 16'h9c28,
// 16'h99f3, 16'h99c9, 16'h9bb4, 16'h9fa7,
// 16'ha58d, 16'had4a, 16'hb6b0, 16'hc19a,
// 16'hcdbd, 16'hdaf1, 16'he8d9, 16'hf743,
// 16'h05d6, 16'h1448, 16'h2259, 16'h2fad,
// 16'h3c14, 16'h473d, 16'h50f5, 16'h590c,
// 16'h5f51, 16'h63ac, 16'h65fe, 16'h6641,
// 16'h6472, 16'h6096, 16'h5acb, 16'h5323,
// 16'h49d1, 16'h3efd, 16'h32e2, 16'h25bf,
// 16'h17db, 16'h0977, 16'hfae7, 16'hec6c,
// 16'hde5b, 16'hd0f4, 16'hc486, 16'hb94b,
// 16'haf7b, 16'ha754, 16'ha0f0, 16'h9c82,
// 16'h9a13, 16'h99b5, 16'h9b6c, 16'h9f2a,
// 16'ha4e2, 16'hac6e, 16'hb5af, 16'hc072,
// 16'hcc79, 16'hd998, 16'he76a, 16'hf5d4,
// 16'h045c, 16'h12dd, 16'h20f7, 16'h2e60,
// 16'h3ae7, 16'h462b, 16'h5011, 16'h5851,
// 16'h5ec5, 16'h6355, 16'h65d9, 16'h6653,
// 16'h64b7, 16'h6112, 16'h5b73, 16'h53fd,
// 16'h4ad1, 16'h4020, 16'h3427, 16'h2719,
// 16'h1945, 16'h0aec, 16'hfc5a, 16'heddc,
// 16'hdfbd, 16'hd240, 16'hc5ba, 16'hba56,
// 16'hb069, 16'ha80d, 16'ha181, 16'h9cda,
// 16'h9a3b, 16'h99a5, 16'h9b2a, 16'h9eb2,
// 16'ha43a, 16'hab98, 16'hb4b1, 16'hbf4d,
// 16'hcb3b, 16'hd83a, 16'he604, 16'hf45d,
// 16'h02ea, 16'h116c, 16'h1f94, 16'h2d14,
// 16'h39b0, 16'h451f, 16'h4f20, 16'h5796,
// 16'h5e33, 16'h62f9, 16'h65af, 16'h6660,
// 16'h64f5, 16'h618a, 16'h5c15, 16'h54d4,
// 16'h4bcb, 16'h4145, 16'h3563, 16'h2874,
// 16'h1aac, 16'h0c61, 16'hfdcf, 16'hef4b,
// 16'he121, 16'hd38f, 16'hc6ef, 16'hbb6a,
// 16'hb156, 16'ha8cd, 16'ha215, 16'h9d3a,
// 16'h9a66, 16'h999d, 16'h9ae9, 16'h9e43,
// 16'ha394, 16'haacb, 16'hb3b1, 16'hbe31,
// 16'hc9f9, 16'hd6e5, 16'he49c, 16'hf2ea,
// 16'h0173, 16'h0ffd, 16'h1e2e, 16'h2bc6,
// 16'h3879, 16'h4409, 16'h4e32, 16'h56d0,
// 16'h5da1, 16'h6294, 16'h6582, 16'h6666,
// 16'h6532, 16'h61f6, 16'h5cbc, 16'h559b,
// 16'h4ccb, 16'h425e, 16'h36a5, 16'h29c6,
// 16'h1c18, 16'h0dce, 16'hff49, 16'hf0bb,
// 16'he284, 16'hd4e5, 16'hc820, 16'hbc89,
// 16'hb240, 16'ha998, 16'ha2aa, 16'h9d9f,
// 16'h9a98, 16'h9999, 16'h9ab0, 16'h9dd6,
// 16'ha2f7, 16'ha9f9, 16'hb2c1, 16'hbd0e,
// 16'hc8c3, 16'hd58b, 16'he339, 16'hf173,
// 16'h2002, 16'h0e8a, 16'h1cc8, 16'h2a75,
// 16'h373e, 16'h42ef, 16'h4d43, 16'h5604,
// 16'h5d0a, 16'h622b, 16'h654d, 16'h6669,
// 16'h6568, 16'h6261, 16'h5d55, 16'h566b,
// 16'h4dba, 16'h437e, 16'h37db, 16'h2b1d,
// 16'h1d7d, 16'h0f41, 16'h20be, 16'hf22b,
// 16'he3ee, 16'hd634, 16'hc960, 16'hbd9d,
// 16'hb33b, 16'haa5f, 16'ha348, 16'h9e08,
// 16'h9acf, 16'h9999, 16'h9a7e, 16'h9d6d,
// 16'ha25e, 16'ha931, 16'hb1ce, 16'hbbf5,
// 16'hc789, 16'hd43a, 16'he1d1, 16'hf004,
// 16'hfe8d, 16'h0d14, 16'h1b66, 16'h291b,
// 16'h3605, 16'h41d3, 16'h4c4b, 16'h5536,
// 16'h5c6e, 16'h61ba, 16'h651a, 16'h6661,
// 16'h659b, 16'h62c4, 16'h5def, 16'h572e,
// 16'h4eb0, 16'h4490, 16'h3916, 16'h2c6e,
// 16'h1ee0, 16'h10b6, 16'h022f, 16'hf3a0,
// 16'he555, 16'hd78a, 16'hca9e, 16'hbebc,
// 16'hb431, 16'hab33, 16'ha3e3, 16'h9e7d,
// 16'h9b06, 16'h99a3, 16'h9a4e, 16'h9d0b,
// 16'ha1c8, 16'ha870, 16'hb0da, 16'hbae5,
// 16'hc64e, 16'hd2ed, 16'he06b, 16'hee96,
// 16'hfd13, 16'h0ba6, 16'h19fa, 16'h27c6,
// 16'h34c6, 16'h40b2, 16'h4b4f, 16'h5468,
// 16'h5bc7, 16'h614b, 16'h64da, 16'h6657,
// 16'h65c8, 16'h6324, 16'h5e80, 16'h57f2,
// 16'h4f99, 16'h45a8, 16'h3a46, 16'h2dc1,
// 16'h2041, 16'h1228, 16'h03a1, 16'hf518,
// 16'he6b9, 16'hd8e7, 16'hcbda, 16'hbfdf,
// 16'hb530, 16'hac04, 16'ha48a, 16'h9ef1,
// 16'h9b46, 16'h99b0, 16'h9a24, 16'h9cae,
// 16'ha139, 16'ha7af, 16'haff1, 16'hb9d1,
// 16'hc51d, 16'hd19e, 16'hdf09, 16'hed25,
// 16'hfb9f, 16'h0a34, 16'h188d, 16'h2670,
// 16'h3381, 16'h3f91, 16'h4a51, 16'h5391,
// 16'h5b1f, 16'h60d6, 16'h6493, 16'h664d,
// 16'h65ea, 16'h6384, 16'h5f08, 16'h58b4,
// 16'h507e, 16'h46ba, 16'h3b79, 16'h2f0b,
// 16'h21a6, 16'h1392, 16'h051c, 16'hf687,
// 16'he827, 16'hda3f, 16'hcd1e, 16'hc104,
// 16'hb62f, 16'hacde, 16'ha533, 16'h9f6b,
// 16'h9b8d, 16'h99c0, 16'h9a02, 16'h9c54,
// 16'ha0af, 16'ha6f3, 16'haf0c, 16'hb8c1,
// 16'hc3f0, 16'hd04e, 16'hddac, 16'hebb4,
// 16'hfa2c, 16'h08be, 16'h1723, 16'h2514,
// 16'h323f, 16'h3e69, 16'h494e, 16'h52b6,
// 16'h5a75, 16'h6057, 16'h644d, 16'h6637,
// 16'h660d, 16'h63d7, 16'h5f95, 16'h5967,
// 16'h5168, 16'h47c3, 16'h3ca7, 16'h3058,
// 16'h2303, 16'h1504, 16'h068d, 16'hf7fd,
// 16'he991, 16'hdb9d, 16'hce62, 16'hc22e,
// 16'hb732, 16'hadba, 16'ha5e4, 16'h9fe7,
// 16'h9bda, 16'h99d7, 16'h99e1, 16'h9c04,
// 16'ha026, 16'ha63f, 16'hae28, 16'hb7b8,
// 16'hc2c1, 16'hcf08, 16'hdc49, 16'hea4b,
// 16'hf8b3, 16'h074c, 16'h15b6, 16'h23b8,
// 16'h30f6, 16'h3d42, 16'h4845, 16'h51d9,
// 16'h59c3, 16'h5fd5, 16'h6402, 16'h6619,
// 16'h662f, 16'h6420, 16'h601f, 16'h5a17,
// 16'h524a, 16'h48ca, 16'h3dd4, 16'h319e,
// 16'h2464, 16'h166e, 16'h0803, 16'hf971,
// 16'heaff, 16'hdcfa, 16'hcfac, 16'hc355,
// 16'hb83f, 16'hae98, 16'ha699, 16'ha06b,
// 16'h9c29, 16'h99f2, 16'h99cb, 16'h9bb2,
// 16'h9faa, 16'ha58a, 16'had4b, 16'hb6b0,
// 16'hc199, 16'hcdbf, 16'hdaef, 16'he8db,
// 16'hf741, 16'h05d6, 16'h1449, 16'h2258,
// 16'h2faf, 16'h3c12, 16'h473d, 16'h50f5,
// 16'h590c, 16'h5f53, 16'h63aa, 16'h65ff,
// 16'h6641, 16'h6470, 16'h609a, 16'h5ac8,
// 16'h5325, 16'h49d0, 16'h3efc, 16'h32e3,
// 16'h25c0, 16'h17d9, 16'h0979, 16'hfae5,
// 16'hec6d, 16'hde5a, 16'hd0f6, 16'hc485,
// 16'hb94a, 16'haf7d, 16'ha752, 16'ha0f1,
// 16'h9c83, 16'h9a10, 16'h99b8, 16'h9b6a,
// 16'h9f2b, 16'ha4e1, 16'hac6e, 16'hb5b0,
// 16'hc070, 16'hcc7d, 16'hd991, 16'he772,
// 16'hf5cc, 16'h0463, 16'h12d9, 16'h20f7,
// 16'h2e63, 16'h3ae3, 16'h462f, 16'h500e,
// 16'h5852, 16'h5ec5, 16'h6356, 16'h65d7,
// 16'h6656, 16'h64b4, 16'h6113, 16'h5b73,
// 16'h53fd, 16'h4ad1, 16'h4022, 16'h3423,
// 16'h271c, 16'h1943, 16'h0aee, 16'hfc59,
// 16'heddc, 16'hdfbc, 16'hd243, 16'hc5b6,
// 16'hba5c, 16'hb062, 16'ha812, 16'ha17d,
// 16'h9cde, 16'h9a39, 16'h99a6, 16'h9b29,
// 16'h9eb1, 16'ha43c, 16'hab97, 16'hb4b3,
// 16'hbf4a, 16'hcb3d, 16'hd838, 16'he608,
// 16'hf459, 16'h02ec, 16'h116b, 16'h1f94,
// 16'h2d15, 16'h39b0, 16'h451d, 16'h4f23,
// 16'h5793, 16'h5e34, 16'h62fa, 16'h65af,
// 16'h665e, 16'h64f9, 16'h6184, 16'h5c1c,
// 16'h54ce, 16'h4bcf, 16'h4142, 16'h3566,
// 16'h2872, 16'h1aae, 16'h0c5e, 16'hfdd2,
// 16'hef49, 16'he122, 16'hd38f, 16'hc6ef,
// 16'hbb6a, 16'hb156, 16'ha8cd, 16'ha214,
// 16'h9d3b, 16'h9a65, 16'h999f, 16'h9ae8,
// 16'h9e42, 16'ha396, 16'haac7, 16'hb3b7,
// 16'hbe2b, 16'hc9fe, 16'hd6e0, 16'he4a1,
// 16'hf2e5, 16'h0178, 16'h0ff8, 16'h1e33,
// 16'h2bc2, 16'h387b, 16'h4408, 16'h4e32,
// 16'h56d2, 16'h5d9e, 16'h6297, 16'h657f,
// 16'h6668, 16'h6532, 16'h61f6, 16'h5cba,
// 16'h559f, 16'h4cc8, 16'h4260, 16'h36a4,
// 16'h29c5, 16'h1c1b, 16'h0dcc, 16'hff4a,
// 16'hf0b9, 16'he287, 16'hd4e2, 16'hc823,
// 16'hbc85, 16'hb243, 16'ha998, 16'ha2a8,
// 16'h9da2, 16'h9a94, 16'h999c, 16'h9ab0,
// 16'h9dd4, 16'ha2f9, 16'ha9f9, 16'hb2bf,
// 16'hbd12, 16'hc8be, 16'hd58f, 16'he336,
// 16'hf176, 16'h2001, 16'h0e89, 16'h1cca,
// 16'h2a72, 16'h3741, 16'h42ee, 16'h4d43,
// 16'h5603, 16'h5d0c, 16'h6227, 16'h6554,
// 16'h6661, 16'h656f, 16'h625b, 16'h5d5a,
// 16'h5667, 16'h4dbe, 16'h437b, 16'h37dc,
// 16'h2b1f, 16'h1d79, 16'h0f46, 16'h20b8,
// 16'hf230, 16'he3eb, 16'hd635, 16'hc960,
// 16'hbd9d, 16'hb33b, 16'haa60, 16'ha345,
// 16'h9e0b, 16'h9acd, 16'h999b, 16'h9a7d,
// 16'h9d6d, 16'ha25d, 16'ha933, 16'hb1cc,
// 16'hbbf6, 16'hc789, 16'hd43a, 16'he1d0,
// 16'hf007, 16'hfe87, 16'h0d1c, 16'h1b5e,
// 16'h2922, 16'h3620, 16'h41d5, 16'h4c4a,
// 16'h5538, 16'h5c6a, 16'h61c0, 16'h6514,
// 16'h6665, 16'h6599, 16'h62c5, 16'h5dee,
// 16'h572f, 16'h4eaf, 16'h4490, 16'h3917,
// 16'h2c6c, 16'h1ee2, 16'h10b4, 16'h0230,
// 16'hf3a1, 16'he552, 16'hd78e, 16'hca9a,
// 16'hbebf, 16'hb430, 16'hab32, 16'ha3e5,
// 16'h9e7b, 16'h9b08, 16'h99a1, 16'h9a50,
// 16'h9d08, 16'ha1cc, 16'ha86c, 16'hb0de,
// 16'hbae1, 16'hc652, 16'hd2ea, 16'he06d,
// 16'hee94, 16'hfd15, 16'h0ba4, 16'h19fd,
// 16'h27c2, 16'h34c9, 16'h40b1, 16'h4b4f,
// 16'h5468, 16'h5bc7, 16'h614c, 16'h64d9,
// 16'h6658, 16'h65c7, 16'h6325, 16'h5e7f,
// 16'h57f4, 16'h4f97, 16'h45a9, 16'h3a47,
// 16'h2dbe, 16'h2045, 16'h1223, 16'h03a7,
// 16'hf512, 16'he6bd, 16'hd8e5, 16'hcbdb,
// 16'hbfe0, 16'hb52c, 16'hac08, 16'ha486,
// 16'h9ef5, 16'h9b44, 16'h99b1, 16'h9a23,
// 16'h9caf, 16'ha136, 16'ha7b3, 16'hafee,
// 16'hb9d3, 16'hc51d, 16'hd19c, 16'hdf0b,
// 16'hed24, 16'hfb9f, 16'h0a34, 16'h188e,
// 16'h266f, 16'h3382, 16'h3f91, 16'h4a4f,
// 16'h5394, 16'h5b1c, 16'h60d9, 16'h6491,
// 16'h664d, 16'h65ec, 16'h6380, 16'h5f0d,
// 16'h58ae, 16'h5084, 16'h46b6, 16'h3b7a,
// 16'h2f0b, 16'h21a5, 16'h1394, 16'h051a,
// 16'hf688, 16'he826, 16'hda40, 16'hcd1e,
// 16'hc103, 16'hb631, 16'hacda, 16'ha538,
// 16'h9f67, 16'h9b8f, 16'h99c0, 16'h9a20,
// 16'h9c57, 16'ha0ac, 16'ha6f5, 16'haf0b,
// 16'hb8c1, 16'hc3f1, 16'hd04d, 16'hddac,
// 16'hebb4, 16'hfa2c, 16'h08bd, 16'h1725,
// 16'h2513, 16'h323e, 16'h3e6b, 16'h494c,
// 16'h52b8, 16'h5a72, 16'h605a, 16'h644c,
// 16'h6635, 16'h6610, 16'h63d5, 16'h5f94,
// 16'h596a, 16'h5164, 16'h47c6, 16'h3ca8,
// 16'h3054, 16'h2306, 16'h1501, 16'h0691,
// 16'hf7fb, 16'he992, 16'hdb9b, 16'hce64,
// 16'hc22c, 16'hb734, 16'hadb8, 16'ha5e5,
// 16'h9fe8, 16'h9bd9, 16'h99d6, 16'h99e3,
// 16'h9c01, 16'ha029, 16'ha63f, 16'hae26,
// 16'hb7bb, 16'hc2be, 16'hcf08, 16'hdc4b,
// 16'hea48, 16'hf8b7, 16'h0749, 16'h15b8,
// 16'h23b5, 16'h30f8, 16'h3d41, 16'h4846,
// 16'h51da, 16'h59c0, 16'h5fd9, 16'h63fe,
// 16'h661d, 16'h662b, 16'h6425, 16'h6019,
// 16'h5a1c, 16'h5247, 16'h48cd, 16'h3dd2,
// 16'h319f, 16'h2461, 16'h1671, 16'h0803,
// 16'hf970, 16'heb20, 16'hdcf8, 16'hcfad,
// 16'hc356, 16'hb83d, 16'hae9a, 16'ha697,
// 16'ha06b, 16'h9c2c, 16'h99ee, 16'h99cf,
// 16'h9baf, 16'h9fa9, 16'ha58d, 16'had48,
// 16'hb6b5, 16'hc194, 16'hcdc2, 16'hdaed,
// 16'he8db, 16'hf744, 16'h05d2, 16'h144e,
// 16'h2253, 16'h2fb2, 16'h3c11, 16'h473d,
// 16'h50f7, 16'h590a, 16'h5f54, 16'h63a8,
// 16'h6602, 16'h663e, 16'h6473, 16'h6097,
// 16'h5aca, 16'h5324, 16'h49d1, 16'h3efb,
// 16'h32e4, 16'h25be, 16'h17dc, 16'h0976,
// 16'hfae7, 16'hec6d, 16'hde5a, 16'hd0f4,
// 16'hc488, 16'hb946, 16'haf81, 16'ha74f,
// 16'ha0f3, 16'h9c81, 16'h9a12, 16'h99b6,
// 16'h9b6c, 16'h9f29, 16'ha4e2, 16'hac6e,
// 16'hb5b0, 16'hc06f, 16'hcc7f, 16'hd98f,
// 16'he773, 16'hf5cd, 16'h0460, 16'h12dc,
// 16'h20f5, 16'h2e64, 16'h3ae2, 16'h4630,
// 16'h500d, 16'h5854, 16'h5ec3, 16'h6356,
// 16'h65d8, 16'h6654, 16'h64b7, 16'h6111,
// 16'h5b74, 16'h53fc, 16'h4ad1, 16'h4022,
// 16'h3424, 16'h271b, 16'h1945, 16'h0aea,
// 16'hfc5e, 16'hedd8, 16'hdfbf, 16'hd240,
// 16'hc5b9, 16'hba59, 16'hb066, 16'ha80e,
// 16'ha180, 16'h9cdc, 16'h9a38, 16'h99a9,
// 16'h9b25, 16'h9eb7, 16'ha436, 16'hab9b,
// 16'hb4af, 16'hbf4e, 16'hcb3b, 16'hd839,
// 16'he607, 16'hf45a, 16'h02eb, 16'h116d,
// 16'h1f91, 16'h2d19, 16'h39ab, 16'h4521,
// 16'h4f21, 16'h5794, 16'h5e35, 16'h62f7,
// 16'h65b0, 16'h665f, 16'h64f9, 16'h6183,
// 16'h5c1e, 16'h54ca, 16'h4bd3, 16'h4140,
// 16'h3566, 16'h2873, 16'h1aad, 16'h0c5e,
// 16'hfdd3, 16'hef48, 16'he123, 16'hd38e,
// 16'hc6ee, 16'hbb6c, 16'hb154, 16'ha8cf,
// 16'ha214, 16'h9d38, 16'h9a69, 16'h999b,
// 16'h9aec, 16'h9e40, 16'ha396, 16'haac9,
// 16'hb3b3, 16'hbe31, 16'hc9f9, 16'hd6e4,
// 16'he49d, 16'hf2e9, 16'h0174, 16'h0ffd,
// 16'h1e2e, 16'h2bc6, 16'h3879, 16'h4407,
// 16'h4e35, 16'h56ce, 16'h5da2, 16'h6293,
// 16'h6583, 16'h6664, 16'h6535, 16'h61f3,
// 16'h5cbc, 16'h559e, 16'h4cc8, 16'h4260,
// 16'h36a2, 16'h29ca, 16'h1c13, 16'h0dd5,
// 16'hff42, 16'hf0c0, 16'he280, 16'hd4e7,
// 16'hc820, 16'hbc88, 16'hb241, 16'ha998,
// 16'ha2a9, 16'h9da0, 16'h9a96, 16'h999b,
// 16'h9aaf, 16'h9dd7, 16'ha2f5, 16'ha9fc,
// 16'hb2be, 16'hbd11, 16'hc8c0, 16'hd58d,
// 16'he337, 16'hf176, 16'h2020, 16'h0e8a,
// 16'h1cca, 16'h2a71, 16'h3742, 16'h42ed,
// 16'h4d44, 16'h5603, 16'h5d0b, 16'h6229,
// 16'h6551, 16'h6665, 16'h656b, 16'h625e,
// 16'h5d59, 16'h5667, 16'h4dbe, 16'h437a,
// 16'h37de, 16'h2b1c, 16'h1d7d, 16'h0f42,
// 16'h20bb, 16'hf22f, 16'he3ea, 16'hd638,
// 16'hc95e, 16'hbd9d, 16'hb33c, 16'haa5e,
// 16'ha349, 16'h9e07, 16'h9ad0, 16'h9998,
// 16'h9a80, 16'h9d6b, 16'ha25f, 16'ha930,
// 16'hb1ce, 16'hbbf7, 16'hc787, 16'hd43b,
// 16'he1d0, 16'hf005, 16'hfe8b, 16'h0d18,
// 16'h1b62, 16'h291e, 16'h3603, 16'h41d3,
// 16'h4c4a, 16'h553a, 16'h5c68, 16'h61c1,
// 16'h6514, 16'h6663, 16'h659b, 16'h62c4,
// 16'h5def, 16'h572f, 16'h4ead, 16'h4494,
// 16'h3912, 16'h2c71, 16'h1ede, 16'h10b7,
// 16'h022e, 16'hf3a2, 16'he552, 16'hd78c,
// 16'hca9e, 16'hbeba, 16'hb434, 16'hab2f,
// 16'ha3e7, 16'h9e79, 16'h9b0a, 16'h999f,
// 16'h9a51, 16'h9d0a, 16'ha1c7, 16'ha872,
// 16'hb0d8, 16'hbae7, 16'hc64e, 16'hd2ec,
// 16'he06b, 16'hee95, 16'hfd17, 16'h0ba2,
// 16'h19fd, 16'h27c3, 16'h34c7, 16'h40b4,
// 16'h4b4d, 16'h546a, 16'h5bc4, 16'h614f,
// 16'h64d7, 16'h6659, 16'h65c7, 16'h6324,
// 16'h5e81, 16'h57f1, 16'h4f9a, 16'h45a7,
// 16'h3a48, 16'h2dbf, 16'h2042, 16'h1226,
// 16'h03a5, 16'hf514, 16'he6bc, 16'hd8e4,
// 16'hcbdd, 16'hbfdd, 16'hb531, 16'hac01,
// 16'ha48f, 16'h9eec, 16'h9b4b, 16'h99ac,
// 16'h9a26, 16'h9cad, 16'ha13a, 16'ha7ad,
// 16'haff4, 16'hb9cf, 16'hc51e, 16'hd19d,
// 16'hdf09, 16'hed26, 16'hfb9f, 16'h0a33,
// 16'h188e, 16'h266f, 16'h3383, 16'h3f8f,
// 16'h4a52, 16'h5390, 16'h5b20, 16'h60d4,
// 16'h6496, 16'h6649, 16'h65f0, 16'h637b,
// 16'h5f11, 16'h58ac, 16'h5085, 16'h46b5,
// 16'h3b7b, 16'h2f0a, 16'h21a7, 16'h1391,
// 16'h051d, 16'hf686, 16'he828, 16'hda3e,
// 16'hcd1f, 16'hc103, 16'hb630, 16'hacdd,
// 16'ha534, 16'h9f6a, 16'h9b8d, 16'h99c1,
// 16'h9a20, 16'h9c57, 16'ha0ab, 16'ha6f6,
// 16'haf0a, 16'hb8c3, 16'hc3ef, 16'hd04e,
// 16'hddac, 16'hebb3, 16'hfa2e, 16'h08bc,
// 16'h1726, 16'h2511, 16'h3240, 16'h3e69,
// 16'h494e, 16'h52b7, 16'h5a72, 16'h605a,
// 16'h644c, 16'h6636, 16'h660e, 16'h63d6,
// 16'h5f95, 16'h5967, 16'h5168, 16'h47c2,
// 16'h3caa, 16'h3055, 16'h2305, 16'h1501,
// 16'h0690, 16'hf7fc, 16'he992, 16'hdb9c,
// 16'hce63, 16'hc22b, 16'hb736, 16'hadb7,
// 16'ha5e6, 16'h9fe6, 16'h9bdb, 16'h99d5,
// 16'h99e4, 16'h9c20, 16'ha02a, 16'ha63c,
// 16'hae2b, 16'hb7b5, 16'hc2c4, 16'hcf03,
// 16'hdc50, 16'hea43, 16'hf8bb, 16'h0746,
// 16'h15b9, 16'h23b6, 16'h30f8, 16'h3d41,
// 16'h4845, 16'h51da, 16'h59c0, 16'h5fda,
// 16'h63fd, 16'h661d, 16'h662b, 16'h6425,
// 16'h601a, 16'h5a1b, 16'h5248, 16'h48cb,
// 16'h3dd4, 16'h319d, 16'h2465, 16'h166d,
// 16'h0805, 16'hf96f, 16'heaff, 16'hdcfc,
// 16'hcfa8, 16'hc35a, 16'hb83b, 16'hae9a,
// 16'ha698, 16'ha06b, 16'h9c29, 16'h99f3,
// 16'h99ca, 16'h9bb3, 16'h9fa8, 16'ha58c,
// 16'had49, 16'hb6b4, 16'hc194, 16'hcdc4,
// 16'hdaea, 16'he8df, 16'hf73f, 16'h05d7,
// 16'h144a, 16'h2256, 16'h2fb0, 16'h3c12,
// 16'h473d, 16'h50f6, 16'h590c, 16'h5f50,
// 16'h63ae, 16'h65fc, 16'h6643, 16'h6470,
// 16'h6098, 16'h5ac9, 16'h5326, 16'h49cf,
// 16'h3efc, 16'h32e4, 16'h25be, 16'h17db,
// 16'h0978, 16'hfae6, 16'hec6c, 16'hde5b,
// 16'hd0f4, 16'hc487, 16'hb949, 16'haf7e,
// 16'ha74f, 16'ha0f5, 16'h9c80, 16'h9a12,
// 16'h99b7, 16'h9b6a, 16'h9f2b, 16'ha4e2,
// 16'hac6d, 16'hb5b1, 16'hc06f, 16'hcc7e,
// 16'hd990, 16'he774, 16'hf5cb, 16'h0462,
// 16'h12da, 16'h20f7, 16'h2e63, 16'h3ae3,
// 16'h462e, 16'h5010, 16'h584f, 16'h5ec9,
// 16'h6352, 16'h65da, 16'h6653, 16'h64b6,
// 16'h6113, 16'h5b72, 16'h53ff, 16'h4ace,
// 16'h4024, 16'h3423, 16'h271b, 16'h1945,
// 16'h0aeb, 16'hfc5c, 16'heddb, 16'hdfbb,
// 16'hd244, 16'hc5b6, 16'hba5a, 16'hb066,
// 16'ha80e, 16'ha180, 16'h9cdc, 16'h9a38,
// 16'h99a9, 16'h9b26, 16'h9eb5, 16'ha438,
// 16'hab99, 16'hb4b2, 16'hbf4c, 16'hcb3a,
// 16'hd83c, 16'he603, 16'hf45f, 16'h02e6,
// 16'h1170, 16'h1f90, 16'h2d18, 16'h39ae,
// 16'h451e, 16'h4f22, 16'h5795, 16'h5e33,
// 16'h62f8, 16'h65b1, 16'h665d, 16'h64fa,
// 16'h6184, 16'h5c1a, 16'h54d0, 16'h4bce,
// 16'h4143, 16'h3564, 16'h2874, 16'h1aad,
// 16'h0c5f, 16'hfdd0, 16'hef4c, 16'he11f,
// 16'hd393, 16'hc6ea, 16'hbb6d, 16'hb155,
// 16'ha8ce, 16'ha214, 16'h9d3b, 16'h9a64,
// 16'h999f, 16'h9ae9, 16'h9e42, 16'ha396,
// 16'haac7, 16'hb3b6, 16'hbe2d, 16'hc9fc,
// 16'hd6e3, 16'he49d, 16'hf2e8, 16'h0175,
// 16'h0ffc, 16'h1e2e, 16'h2bc8, 16'h3875,
// 16'h440c, 16'h4e30, 16'h56d2, 16'h5da0,
// 16'h6294, 16'h6583, 16'h6664, 16'h6534,
// 16'h61f5, 16'h5cba, 16'h55a0, 16'h4cc6,
// 16'h4262, 16'h36a1, 16'h29ca, 16'h1c15,
// 16'h0dd0, 16'hff49, 16'hf0b8, 16'he289,
// 16'hd4e0, 16'hc824, 16'hbc86, 16'hb241,
// 16'ha999, 16'ha2a8, 16'h9da1, 16'h9a96,
// 16'h999a, 16'h9aaf, 16'h9dd8, 16'ha2f4,
// 16'ha9fe, 16'hb2bb, 16'hbd13, 16'hc8bf,
// 16'hd58e, 16'he338, 16'hf174, 16'h2002,
// 16'h0e87, 16'h1ccd, 16'h2a6f, 16'h3744,
// 16'h42ec, 16'h4d43, 16'h5605, 16'h5d07,
// 16'h622e, 16'h654d, 16'h6667, 16'h656b,
// 16'h625d, 16'h5d5a, 16'h5665, 16'h4dc1,
// 16'h4378, 16'h37df, 16'h2b1c, 16'h1d7b,
// 16'h0f45, 16'h20b9, 16'hf230, 16'he3e9,
// 16'hd639, 16'hc95c, 16'hbda0, 16'hb339,
// 16'haa61, 16'ha344, 16'h9e0e, 16'h9ac9,
// 16'h999e, 16'h9a7b, 16'h9d6e, 16'ha25e,
// 16'ha932, 16'hb1cb, 16'hbbf8, 16'hc788,
// 16'hd43a, 16'he1d1, 16'hf004, 16'hfe8c,
// 16'h0d16, 16'h1b64, 16'h291c, 16'h3606,
// 16'h41d0, 16'h4c4d, 16'h5537, 16'h5c6b,
// 16'h61bf, 16'h6514, 16'h6665, 16'h6598,
// 16'h62c8, 16'h5dea, 16'h5733, 16'h4eab,
// 16'h4494, 16'h3914, 16'h2c6d, 16'h1ee2,
// 16'h10b4, 16'h0230, 16'hf3a1, 16'he552,
// 16'hd78e, 16'hca9a, 16'hbebf, 16'hb42f,
// 16'hab33, 16'ha3e5, 16'h9e7b, 16'h9b07,
// 16'h99a3, 16'h9a4d, 16'h9d0d, 16'ha1c6,
// 16'ha871, 16'hb0da, 16'hbae4, 16'hc651,
// 16'hd2ea, 16'he06c, 16'hee96, 16'hfd13,
// 16'h0ba7, 16'h19f9, 16'h27c6, 16'h34c7,
// 16'h40b1, 16'h4b50, 16'h5467, 16'h5bc8,
// 16'h614b, 16'h64da, 16'h6656, 16'h65c9,
// 16'h6324, 16'h5e80, 16'h57f1, 16'h4f9c,
// 16'h45a3, 16'h3a4d, 16'h2db9, 16'h2048,
// 16'h1222, 16'h03a7, 16'hf513, 16'he6bc,
// 16'hd8e5, 16'hcbdc, 16'hbfdf, 16'hb52e,
// 16'hac05, 16'ha48b, 16'h9eef, 16'h9b4a,
// 16'h99ac, 16'h9a26, 16'h9cae, 16'ha138,
// 16'ha7af, 16'haff3, 16'hb9cd, 16'hc523,
// 16'hd197, 16'hdf0e, 16'hed22, 16'hfba1,
// 16'h0a32, 16'h188f, 16'h266d, 16'h3385,
// 16'h3f8e, 16'h4a52, 16'h5390, 16'h5b1f,
// 16'h60d6, 16'h6495, 16'h6649, 16'h65ef,
// 16'h637c, 16'h5f13, 16'h58a8, 16'h508a,
// 16'h46b0, 16'h3b7f, 16'h2f08, 16'h21a7,
// 16'h1393, 16'h051a, 16'hf689, 16'he825,
// 16'hda40, 16'hcd1e, 16'hc103, 16'hb631,
// 16'hacda, 16'ha538, 16'h9f67, 16'h9b90,
// 16'h99be, 16'h9a02, 16'h9c54, 16'ha0af,
// 16'ha6f5, 16'haf08, 16'hb8c7, 16'hc3e9,
// 16'hd055, 16'hdda6, 16'hebb8, 16'hfa2a,
// 16'h08be, 16'h1725, 16'h2512, 16'h3240,
// 16'h3e68, 16'h494f, 16'h52b6, 16'h5a74,
// 16'h6058, 16'h644d, 16'h6635, 16'h6611,
// 16'h63d2, 16'h5f9a, 16'h5962, 16'h516c,
// 16'h47bf, 16'h3cac, 16'h3053, 16'h2307,
// 16'h1501, 16'h068e, 16'hf7ff, 16'he98d,
// 16'hdba1, 16'hce60, 16'hc22d, 16'hb735,
// 16'hadb6, 16'ha5e7, 16'h9fe6, 16'h9bda,
// 16'h99d7, 16'h99e0, 16'h9c05, 16'ha026,
// 16'ha63f, 16'hae28, 16'hb7b8, 16'hc2c0,
// 16'hcf09, 16'hdc49, 16'hea4a, 16'hf8b4,
// 16'h074c, 16'h15b5, 16'h23b9, 16'h30f6,
// 16'h3d41, 16'h4846, 16'h51d9, 16'h59c2,
// 16'h5fd7, 16'h63ff, 16'h661d, 16'h662a,
// 16'h6426, 16'h6019, 16'h5a1b, 16'h5248,
// 16'h48cc, 16'h3dd3, 16'h319e, 16'h2463,
// 16'h166f, 16'h0804, 16'hf970, 16'heb20,
// 16'hdcf8, 16'hcfae, 16'hc354, 16'hb841,
// 16'hae94, 16'ha69d, 16'ha067, 16'h9c2d,
// 16'h99f1, 16'h99c9, 16'h9bb5, 16'h9fa5,
// 16'ha58f, 16'had49, 16'hb6b0, 16'hc19a,
// 16'hcdbd, 16'hdaf1, 16'he8d9, 16'hf743,
// 16'h05d5, 16'h144a, 16'h2257, 16'h2faf,
// 16'h3c12, 16'h473e, 16'h50f5, 16'h590c,
// 16'h5f51, 16'h63ad, 16'h65fd, 16'h6642,
// 16'h646f, 16'h609b, 16'h5ac6, 16'h5329,
// 16'h49cb, 16'h3f20, 16'h32e1, 16'h25bf,
// 16'h17dc, 16'h0976, 16'hfae8, 16'hec6b,
// 16'hde5a, 16'hd0f6, 16'hc486, 16'hb949,
// 16'haf7e, 16'ha750, 16'ha0f4, 16'h9c80,
// 16'h9a12, 16'h99b8, 16'h9b68, 16'h9f2e,
// 16'ha4de, 16'hac70, 16'hb5b0, 16'hc06e,
// 16'hcc7f, 16'hd991, 16'he771, 16'hf5ce,
// 16'h0460, 16'h12db, 16'h20f7, 16'h2e63,
// 16'h3ae2, 16'h4630, 16'h500e, 16'h5850,
// 16'h5ec9, 16'h6350, 16'h65de, 16'h6650,
// 16'h64b7, 16'h6113, 16'h5b72, 16'h53fe,
// 16'h4ad0, 16'h4021, 16'h3426, 16'h2719,
// 16'h1946, 16'h0aea, 16'hfc5c, 16'heddb,
// 16'hdfbc, 16'hd243, 16'hc5b6, 16'hba5b,
// 16'hb064, 16'ha811, 16'ha17e, 16'h9cdd,
// 16'h9a37, 16'h99aa, 16'h9b25, 16'h9eb6,
// 16'ha438, 16'hab98, 16'hb4b2, 16'hbf4b,
// 16'hcb3e, 16'hd836, 16'he609, 16'hf458,
// 16'h02ed, 16'h116b, 16'h1f93, 16'h2d17,
// 16'h39ad, 16'h451f, 16'h4f23, 16'h5791,
// 16'h5e39, 16'h62f3, 16'h65b4, 16'h665d,
// 16'h64f7, 16'h6188, 16'h5c17, 16'h54d2,
// 16'h4bce, 16'h4142, 16'h3565, 16'h2873,
// 16'h1aad, 16'h0c60, 16'hfdcf, 16'hef4d,
// 16'he11e, 16'hd392, 16'hc6ec, 16'hbb6d,
// 16'hb152, 16'ha8d2, 16'ha211, 16'h9d3c,
// 16'h9a65, 16'h999d, 16'h9aea, 16'h9e43,
// 16'ha394, 16'haac9, 16'hb3b4, 16'hbe2f,
// 16'hc9fb, 16'hd6e3, 16'he49e, 16'hf2e7,
// 16'h0176, 16'h0ffc, 16'h1e2f, 16'h2bc4,
// 16'h387c, 16'h4403, 16'h4e3a, 16'h56ca,
// 16'h5da5, 16'h6291, 16'h6584, 16'h6664,
// 16'h6534, 16'h61f6, 16'h5cb9, 16'h55a0,
// 16'h4cc7, 16'h4260, 16'h36a4, 16'h29c6,
// 16'h1c18, 16'h0dd0, 16'hff46, 16'hf0bd,
// 16'he283, 16'hd4e4, 16'hc824, 16'hbc83,
// 16'hb245, 16'ha995, 16'ha2ab, 16'h9da0,
// 16'h9a96, 16'h999a, 16'h9aaf, 16'h9dd8,
// 16'ha2f5, 16'ha9fc, 16'hb2bd, 16'hbd11,
// 16'hc8c1, 16'hd58e, 16'he335, 16'hf178,
// 16'hfffc, 16'h0e8f, 16'h1cc5, 16'h2a77,
// 16'h373d, 16'h42ef, 16'h4d43, 16'h5603,
// 16'h5d0d, 16'h6227, 16'h6552, 16'h6665,
// 16'h6569, 16'h6263, 16'h5d51, 16'h5670,
// 16'h4db6, 16'h4381, 16'h37d9, 16'h2b1e,
// 16'h1d7c, 16'h0f43, 16'h20bb, 16'hf22e,
// 16'he3ea, 16'hd639, 16'hc95c, 16'hbda1,
// 16'hb337, 16'haa61, 16'ha347, 16'h9e0a,
// 16'h9acd, 16'h999b, 16'h9a7c, 16'h9d6f,
// 16'ha25b, 16'ha936, 16'hb1c8, 16'hbbf9,
// 16'hc789, 16'hd437, 16'he1d4, 16'hf003,
// 16'hfe8b, 16'h0d19, 16'h1b60, 16'h2920,
// 16'h3602, 16'h41d3, 16'h4c4c, 16'h5537,
// 16'h5c6b, 16'h61bf, 16'h6514, 16'h6664,
// 16'h659b, 16'h62c4, 16'h5def, 16'h572e,
// 16'h4eae, 16'h4493, 16'h3914, 16'h2c6f,
// 16'h1ee0, 16'h10b4, 16'h0231, 16'hf3a1,
// 16'he551, 16'hd790, 16'hca98, 16'hbec0,
// 16'hb430, 16'hab31, 16'ha3e6, 16'h9e7b,
// 16'h9b08, 16'h99a1, 16'h9a4f, 16'h9d0a,
// 16'ha1ca, 16'ha86e, 16'hb0db, 16'hbae5,
// 16'hc64e, 16'hd2ed, 16'he06b, 16'hee94,
// 16'hfd16, 16'h0ba5, 16'h19f9, 16'h27c8,
// 16'h34c3, 16'h40b4, 16'h4b51, 16'h5464,
// 16'h5bcb, 16'h6148, 16'h64db, 16'h6658,
// 16'h65c7, 16'h6325, 16'h5e7f, 16'h57f3,
// 16'h4f97, 16'h45ab, 16'h3a44, 16'h2dc2,
// 16'h2041, 16'h1226, 16'h03a4, 16'hf515,
// 16'he6bc, 16'hd8e4, 16'hcbdd, 16'hbfdd,
// 16'hb52f, 16'hac06, 16'ha489, 16'h9ef1,
// 16'h9b47, 16'h99af, 16'h9a25, 16'h9cad,
// 16'ha13a, 16'ha7ae, 16'haff1, 16'hb9d2,
// 16'hc51d, 16'hd19c, 16'hdf0d, 16'hed20,
// 16'hfba4, 16'h0a2f, 16'h1892, 16'h266c,
// 16'h3385, 16'h3f8e, 16'h4a51, 16'h5392,
// 16'h5b1f, 16'h60d5, 16'h6495, 16'h6649,
// 16'h65ee, 16'h6381, 16'h5f0b, 16'h58b0,
// 16'h5082, 16'h46b7, 16'h3b7a, 16'h2f0b,
// 16'h21a5, 16'h1394, 16'h051b, 16'hf686,
// 16'he828, 16'hda3e, 16'hcd1f, 16'hc104,
// 16'hb62f, 16'hacdd, 16'ha534, 16'h9f6a,
// 16'h9b8e, 16'h99c0, 16'h9a01, 16'h9c55,
// 16'ha0ad, 16'ha6f6, 16'haf09, 16'hb8c5,
// 16'hc3eb, 16'hd052, 16'hdda9, 16'hebb6,
// 16'hfa2b, 16'h08be, 16'h1724, 16'h2513,
// 16'h323f, 16'h3e69, 16'h494f, 16'h52b6,
// 16'h5a72, 16'h605c, 16'h6448, 16'h663b,
// 16'h660a, 16'h63d8, 16'h5f94, 16'h5968,
// 16'h5167, 16'h47c3, 16'h3ca8, 16'h3057,
// 16'h2302, 16'h1505, 16'h068d, 16'hf7fe,
// 16'he990, 16'hdb9e, 16'hce60, 16'hc230,
// 16'hb731, 16'hadbb, 16'ha5e3, 16'h9fe8,
// 16'h9bda, 16'h99d5, 16'h99e4, 16'h9c02,
// 16'ha026, 16'ha641, 16'hae25, 16'hb7bb,
// 16'hc2bf, 16'hcf09, 16'hdc48, 16'hea4a,
// 16'hf8b6, 16'h0749, 16'h15ba, 16'h23b2,
// 16'h30fb, 16'h3d3f, 16'h4847, 16'h51d9,
// 16'h59c0, 16'h5fda, 16'h63fc, 16'h6620,
// 16'h6626, 16'h642a, 16'h6016, 16'h5a1c,
// 16'h524a, 16'h48c7, 16'h3dda, 16'h3196,
// 16'h246a, 16'h166b, 16'h0805, 16'hf971,
// 16'heafd, 16'hdcfc, 16'hcfab, 16'hc356,
// 16'hb83e, 16'hae98, 16'ha699, 16'ha06b,
// 16'h9c2a, 16'h99f2, 16'h99c9, 16'h9bb5,
// 16'h9fa5, 16'ha590, 16'had46, 16'hb6b4,
// 16'hc197, 16'hcdbf, 16'hdaef, 16'he8dc,
// 16'hf740, 16'h05d8, 16'h1448, 16'h2257,
// 16'h2fb0, 16'h3c13, 16'h473b, 16'h50f8,
// 16'h5909, 16'h5f54, 16'h63aa, 16'h6620,
// 16'h663e, 16'h6474, 16'h6096, 16'h5acb,
// 16'h5324, 16'h49d0, 16'h3efc, 16'h32e4,
// 16'h25bd, 16'h17dd, 16'h0976, 16'hfae8,
// 16'hec6a, 16'hde5c, 16'hd0f4, 16'hc486,
// 16'hb94a, 16'haf7c, 16'ha753, 16'ha0f1,
// 16'h9c81, 16'h9a13, 16'h99b5, 16'h9b6c,
// 16'h9f2b, 16'ha4df, 16'hac71, 16'hb5ae,
// 16'hc071, 16'hcc7d, 16'hd991, 16'he771,
// 16'hf5cf, 16'h045e, 16'h12df, 16'h20f2,
// 16'h2e66, 16'h3ae2, 16'h462f, 16'h500e,
// 16'h5852, 16'h5ec6, 16'h6353, 16'h65dd,
// 16'h664e, 16'h64bb, 16'h610e, 16'h5b77,
// 16'h53fa, 16'h4ad3, 16'h401f, 16'h3427,
// 16'h2719, 16'h1946, 16'h0aea, 16'hfc5c,
// 16'heddb, 16'hdfbc, 16'hd243, 16'hc5b6,
// 16'hba5b, 16'hb064, 16'ha811, 16'ha17e,
// 16'h9cdd, 16'h9a37, 16'h99aa, 16'h9b26,
// 16'h9eb5, 16'ha438, 16'hab98, 16'hb4b3,
// 16'hbf4a, 16'hcb3f, 16'hd834, 16'he60c,
// 16'hf456, 16'h02ee, 16'h1169, 16'h1f97,
// 16'h2d12, 16'h39b3, 16'h4519, 16'h4f27,
// 16'h5790, 16'h5e38, 16'h62f5, 16'h65b1,
// 16'h665f, 16'h64f8, 16'h6185, 16'h5c1a,
// 16'h54cf, 16'h4bcf, 16'h4143, 16'h3564,
// 16'h2873, 16'h1aae, 16'h0c5e, 16'hfdd1,
// 16'hef4b, 16'he11f, 16'hd393, 16'hc6ea,
// 16'hbb6f, 16'hb151, 16'ha8d1, 16'ha212,
// 16'h9d3c, 16'h9a65, 16'h999e, 16'h9ae9,
// 16'h9e42, 16'ha395, 16'haac9, 16'hb3b4,
// 16'hbe2f, 16'hc9fb, 16'hd6e2, 16'he49f,
// 16'hf2e6, 16'h0178, 16'h0ffa, 16'h1e2f,
// 16'h2bc6, 16'h3879, 16'h4407, 16'h4e36,
// 16'h56cc, 16'h5da4, 16'h6292, 16'h6583,
// 16'h6665, 16'h6533, 16'h61f6, 16'h5cba,
// 16'h559e, 16'h4cc9, 16'h425f, 16'h36a4,
// 16'h29c7, 16'h1c16, 16'h0dd2, 16'hff45,
// 16'hf0bd, 16'he284, 16'hd4e2, 16'hc826,
// 16'hbc82, 16'hb245, 16'ha996, 16'ha2aa,
// 16'h9d9f, 16'h9a99, 16'h9996, 16'h9ab4,
// 16'h9dd3, 16'ha2f8, 16'ha9fa, 16'hb2bf,
// 16'hbd11, 16'hc8bf, 16'hd590, 16'he334,
// 16'hf178, 16'hfffe, 16'h0e8b, 16'h1cca,
// 16'h2a72, 16'h3740, 16'h42ee, 16'h4d43,
// 16'h5605, 16'h5d08, 16'h622c, 16'h654e,
// 16'h6667, 16'h656b, 16'h625d, 16'h5d59,
// 16'h5667, 16'h4dbe, 16'h437b, 16'h37dc,
// 16'h2b1e, 16'h1d7b, 16'h0f43, 16'h20bc,
// 16'hf22d, 16'he3ec, 16'hd636, 16'hc95f,
// 16'hbd9d, 16'hb33b, 16'haa60, 16'ha346,
// 16'h9e0b, 16'h9acc, 16'h999b, 16'h9a7d,
// 16'h9d6e, 16'ha25d, 16'ha932, 16'hb1cd,
// 16'hbbf5, 16'hc78b, 16'hd437, 16'he1d3,
// 16'hf004, 16'hfe89, 16'h0d1c, 16'h1b5d,
// 16'h2923, 16'h35ff, 16'h41d6, 16'h4c49,
// 16'h5539, 16'h5c6b, 16'h61bd, 16'h6517,
// 16'h6662, 16'h659c, 16'h62c3, 16'h5df0,
// 16'h572c, 16'h4eb1, 16'h4490, 16'h3917,
// 16'h2c6c, 16'h1ee2, 16'h10b3, 16'h0230,
// 16'hf3a3, 16'he551, 16'hd78d, 16'hca9c,
// 16'hbebc, 16'hb434, 16'hab2e, 16'ha3e8,
// 16'h9e79, 16'h9b0a, 16'h999f, 16'h9a51,
// 16'h9d09, 16'ha1cb, 16'ha86c, 16'hb0de,
// 16'hbae1, 16'hc652, 16'hd2eb, 16'he06b,
// 16'hee96, 16'hfd14, 16'h0ba5, 16'h19fa,
// 16'h27c7, 16'h34c4, 16'h40b4, 16'h4b4f,
// 16'h5466, 16'h5bc9, 16'h614b, 16'h64d9,
// 16'h6658, 16'h65c7, 16'h6324, 16'h5e82,
// 16'h57ef, 16'h4f9d, 16'h45a2, 16'h3a4e,
// 16'h2db9, 16'h2048, 16'h1221, 16'h03a7,
// 16'hf514, 16'he6bb, 16'hd8e7, 16'hcbd9,
// 16'hbfe0, 16'hb52e, 16'hac05, 16'ha48b,
// 16'h9eef, 16'h9b49, 16'h99ad, 16'h9a27,
// 16'h9cab, 16'ha13b, 16'ha7ad, 16'haff3,
// 16'hb9d0, 16'hc51f, 16'hd19a, 16'hdf0d,
// 16'hed21, 16'hfba3, 16'h0a31, 16'h188f,
// 16'h266e, 16'h3384, 16'h3f8f, 16'h4a51,
// 16'h5392, 16'h5b1d, 16'h60d8, 16'h6493,
// 16'h664b, 16'h65ed, 16'h6380, 16'h5f0c,
// 16'h58b1, 16'h5080, 16'h46b9, 16'h3b79,
// 16'h2f0a, 16'h21a8, 16'h1390, 16'h051e,
// 16'hf685, 16'he828, 16'hda3e, 16'hcd20,
// 16'hc101, 16'hb633, 16'hacd8, 16'ha539,
// 16'h9f67, 16'h9b8f, 16'h99c0, 16'h9a20,
// 16'h9c56, 16'ha0ad, 16'ha6f6, 16'haf08,
// 16'hb8c5, 16'hc3ed, 16'hd050, 16'hddab,
// 16'hebb4, 16'hfa2c, 16'h08bf, 16'h1721,
// 16'h2516, 16'h323d, 16'h3e6b, 16'h494d,
// 16'h52b7, 16'h5a72, 16'h605b, 16'h644a,
// 16'h6638, 16'h660e, 16'h63d5, 16'h5f96,
// 16'h5967, 16'h5168, 16'h47c2, 16'h3caa,
// 16'h3053, 16'h2308, 16'h1520, 16'h0690,
// 16'hf7fb, 16'he993, 16'hdb9b, 16'hce64,
// 16'hc22b, 16'hb735, 16'hadb8, 16'ha5e4,
// 16'h9fe9, 16'h9bd8, 16'h99d8, 16'h99e1,
// 16'h9c02, 16'ha028, 16'ha63f, 16'hae28,
// 16'hb7b8, 16'hc2c1, 16'hcf06, 16'hdc4b,
// 16'hea4a, 16'hf8b4, 16'h074c, 16'h15b5,
// 16'h23b7, 16'h30f9, 16'h3d3f, 16'h4848,
// 16'h51d7, 16'h59c2, 16'h5fd9, 16'h63fd,
// 16'h661e, 16'h6629, 16'h6427, 16'h6019,
// 16'h5a1a, 16'h524a, 16'h48c8, 16'h3dd8,
// 16'h319b, 16'h2463, 16'h1670, 16'h0803,
// 16'hf970, 16'heb01, 16'hdcf8, 16'hcfac,
// 16'hc357, 16'hb83d, 16'hae98, 16'ha69b,
// 16'ha068, 16'h9c2c, 16'h99f2, 16'h99c8,
// 16'h9bb6, 16'h9fa6, 16'ha58c, 16'had4c,
// 16'hb6ae, 16'hc19b, 16'hcdbd, 16'hdaf1,
// 16'he8d9, 16'hf743, 16'h05d5, 16'h1449,
// 16'h2259, 16'h2fad, 16'h3c14, 16'h473c,
// 16'h50f7, 16'h590a, 16'h5f54, 16'h63a8,
// 16'h6602, 16'h663e, 16'h6473, 16'h6097,
// 16'h5ac9, 16'h5327, 16'h49cc, 16'h3f01,
// 16'h32de, 16'h25c3, 16'h17d9, 16'h0977,
// 16'hfae8, 16'hec6a, 16'hde5c, 16'hd0f5,
// 16'hc486, 16'hb949, 16'haf7d, 16'ha751,
// 16'ha0f4, 16'h9c80, 16'h9a13, 16'h99b6,
// 16'h9b6a, 16'h9f2d, 16'ha4de, 16'hac72,
// 16'hb5ac, 16'hc074, 16'hcc79, 16'hd995,
// 16'he76f, 16'hf5ce, 16'h0461, 16'h12da,
// 16'h20f7, 16'h2e63, 16'h3ae3, 16'h462f,
// 16'h500e, 16'h5852, 16'h5ec5, 16'h6355,
// 16'h65da, 16'h6652, 16'h64b8, 16'h610f,
// 16'h5b77, 16'h53fa, 16'h4ad2, 16'h4021,
// 16'h3425, 16'h271b, 16'h1943, 16'h0aed,
// 16'hfc5a, 16'heddd, 16'hdfbb, 16'hd242,
// 16'hc5b7, 16'hba5a, 16'hb066, 16'ha80f,
// 16'ha17f, 16'h9cdc, 16'h9a39, 16'h99a7,
// 16'h9b28, 16'h9eb4, 16'ha438, 16'hab9b,
// 16'hb4ad, 16'hbf50, 16'hcb3a, 16'hd839,
// 16'he608, 16'hf458, 16'h02ec, 16'h116d,
// 16'h1f91, 16'h2d19, 16'h39ac, 16'h451f,
// 16'h4f23, 16'h5792, 16'h5e37, 16'h62f5,
// 16'h65b3, 16'h665c, 16'h64fa, 16'h6185,
// 16'h5c19, 16'h54d1, 16'h4bcd, 16'h4144,
// 16'h3565, 16'h2871, 16'h1aaf, 16'h0c5f,
// 16'hfdd0, 16'hef4c, 16'he11f, 16'hd391,
// 16'hc6ed, 16'hbb6c, 16'hb155, 16'ha8ce,
// 16'ha214, 16'h9d39, 16'h9a68, 16'h999c,
// 16'h9aeb, 16'h9e40, 16'ha396, 16'haac9,
// 16'hb3b4, 16'hbe2e, 16'hc9fc, 16'hd6e2,
// 16'he49f, 16'hf2e7, 16'h0176, 16'h0ffa,
// 16'h1e31, 16'h2bc5, 16'h3877, 16'h440b,
// 16'h4e32, 16'h56cf, 16'h5da3, 16'h6291,
// 16'h6584, 16'h6665, 16'h6533, 16'h61f6,
// 16'h5cba, 16'h559f, 16'h4cc7, 16'h4260,
// 16'h36a5, 16'h29c5, 16'h1c1a, 16'h0dcd,
// 16'hff48, 16'hf0bc, 16'he284, 16'hd4e4,
// 16'hc823, 16'hbc83, 16'hb246, 16'ha995,
// 16'ha2ab, 16'h9d9e, 16'h9a99, 16'h9997,
// 16'h9ab4, 16'h9dd2, 16'ha2fa, 16'ha9f8,
// 16'hb2c0, 16'hbd10, 16'hc8c1, 16'hd58d,
// 16'he336, 16'hf177, 16'hfffe, 16'h0e8d,
// 16'h1cc7, 16'h2a73, 16'h3740, 16'h42ef,
// 16'h4d41, 16'h5608, 16'h5d05, 16'h622e,
// 16'h654d, 16'h6667, 16'h656b, 16'h625d,
// 16'h5d5a, 16'h5665, 16'h4dc1, 16'h4377,
// 16'h37e0, 16'h2b1b, 16'h1d7d, 16'h0f42,
// 16'h20bd, 16'hf22b, 16'he3ee, 16'hd635,
// 16'hc95e, 16'hbda0, 16'hb338, 16'haa61,
// 16'ha347, 16'h9e08, 16'h9acf, 16'h999a,
// 16'h9a7d, 16'h9d6e, 16'ha25c, 16'ha934,
// 16'hb1cb, 16'hbbf7, 16'hc789, 16'hd438,
// 16'he1d4, 16'hf002, 16'hfe8c, 16'h0d17,
// 16'h1b63, 16'h291e, 16'h3603, 16'h41d3,
// 16'h4c4a, 16'h5539, 16'h5c6a, 16'h61bf,
// 16'h6516, 16'h6661, 16'h659d, 16'h62c3,
// 16'h5def, 16'h572f, 16'h4ead, 16'h4493,
// 16'h3915, 16'h2c6e, 16'h1ee0, 16'h10b5,
// 16'h022f, 16'hf3a3, 16'he550, 16'hd790,
// 16'hca98, 16'hbec0, 16'hb430, 16'hab32,
// 16'ha3e5, 16'h9e7b, 16'h9b07, 16'h99a3,
// 16'h9a4e, 16'h9d0a, 16'ha1ca, 16'ha86d,
// 16'hb0de, 16'hbae0, 16'hc654, 16'hd2e8,
// 16'he06f, 16'hee92, 16'hfd16, 16'h0ba4,
// 16'h19fd, 16'h27c3, 16'h34c7, 16'h40b2,
// 16'h4b50, 16'h5466, 16'h5bc9, 16'h614a,
// 16'h64db, 16'h6657, 16'h65c7, 16'h6324,
// 16'h5e82, 16'h57f0, 16'h4f9b, 16'h45a6,
// 16'h3a48, 16'h2dbf, 16'h2044, 16'h1223,
// 16'h03a7, 16'hf512, 16'he6be, 16'hd8e4,
// 16'hcbdb, 16'hbfe0, 16'hb52e, 16'hac04,
// 16'ha48c, 16'h9eee, 16'h9b4a, 16'h99ae,
// 16'h9a24, 16'h9cae, 16'ha138, 16'ha7b0,
// 16'haff1, 16'hb9d1, 16'hc51d, 16'hd19e,
// 16'hdf07, 16'hed28, 16'hfb9c, 16'h0a36,
// 16'h188d, 16'h266f, 16'h3382, 16'h3f91,
// 16'h4a4f, 16'h5393, 16'h5b1e, 16'h60d5,
// 16'h6497, 16'h6647, 16'h65f1, 16'h637b,
// 16'h5f11, 16'h58ac, 16'h5085, 16'h46b6,
// 16'h3b79, 16'h2f0c, 16'h21a5, 16'h1393,
// 16'h051c, 16'hf686, 16'he827, 16'hda3f,
// 16'hcd1f, 16'hc103, 16'hb62f, 16'hacdd,
// 16'ha535, 16'h9f6a, 16'h9b8d, 16'h99c0,
// 16'h9a01, 16'h9c55, 16'ha0af, 16'ha6f2,
// 16'haf0e, 16'hb8bf, 16'hc3f1, 16'hd04e,
// 16'hddaa, 16'hebb7, 16'hfa2a, 16'h08be,
// 16'h1725, 16'h2512, 16'h323f, 16'h3e6a,
// 16'h494d, 16'h52b8, 16'h5a72, 16'h605a,
// 16'h644a, 16'h6639, 16'h660c, 16'h63d7,
// 16'h5f95, 16'h5968, 16'h5166, 16'h47c4,
// 16'h3ca8, 16'h3056, 16'h2306, 16'h1501,
// 16'h068e, 16'hf7ff, 16'he98e, 16'hdba0,
// 16'hce60, 16'hc22e, 16'hb734, 16'hadb7,
// 16'ha5e7, 16'h9fe5, 16'h9bdb, 16'h99d7,
// 16'h99e0, 16'h9c05, 16'ha025, 16'ha640,
// 16'hae28, 16'hb7b7, 16'hc2c3, 16'hcf05,
// 16'hdc4c, 16'hea48, 16'hf8b6, 16'h074b,
// 16'h15b5, 16'h23b9, 16'h30f5, 16'h3d43,
// 16'h4845, 16'h51d9, 16'h59c2, 16'h5fd7,
// 16'h63ff, 16'h661c, 16'h662c, 16'h6424,
// 16'h601b, 16'h5a19, 16'h5249, 16'h48cc,
// 16'h3dd2, 16'h31a1, 16'h245f, 16'h1672,
// 16'h0802, 16'hf971, 16'heaff, 16'hdcfa,
// 16'hcfab, 16'hc358, 16'hb83c, 16'hae99,
// 16'ha698, 16'ha06c, 16'h9c29, 16'h99f4,
// 16'h99c7, 16'h9bb6, 16'h9fa6, 16'ha58d,
// 16'had4a, 16'hb6b2, 16'hc196, 16'hcdc2,
// 16'hdaec, 16'he8dd, 16'hf741, 16'h05d5,
// 16'h144c, 16'h2254, 16'h2fb2, 16'h3c10,
// 16'h473d, 16'h50f8, 16'h5909, 16'h5f55,
// 16'h63a7, 16'h6602, 16'h663e, 16'h6474,
// 16'h6096, 16'h5aca, 16'h5324, 16'h49d1,
// 16'h3efb, 16'h32e4, 16'h25bf, 16'h17da,
// 16'h0978, 16'hfae6, 16'hec6c, 16'hde5b,
// 16'hd0f5, 16'hc485, 16'hb94b, 16'haf7c,
// 16'ha751, 16'ha0f4, 16'h9c7f, 16'h9a15,
// 16'h99b4, 16'h9b6c, 16'h9f2a, 16'ha4e1,
// 16'hac70, 16'hb5ae, 16'hc072, 16'hcc7b,
// 16'hd993, 16'he770, 16'hf5cf, 16'h045e,
// 16'h12df, 16'h20f3, 16'h2e65, 16'h3ae2,
// 16'h462f, 16'h500e, 16'h5854, 16'h5ec2,
// 16'h6358, 16'h65d6, 16'h6657, 16'h64b2,
// 16'h6116, 16'h5b70, 16'h53ff, 16'h4ad0,
// 16'h4021, 16'h3426, 16'h2719, 16'h1946,
// 16'h0aea, 16'hfc5c, 16'heddc, 16'hdfba,
// 16'hd245, 16'hc5b5, 16'hba5a, 16'hb066,
// 16'ha80f, 16'ha180, 16'h9cdb, 16'h9a39,
// 16'h99a7, 16'h9b28, 16'h9eb5, 16'ha437,
// 16'hab9a, 16'hb4b0, 16'hbf4d, 16'hcb3c,
// 16'hd837, 16'he60a, 16'hf457, 16'h02ee,
// 16'h1169, 16'h1f95, 16'h2d15, 16'h39b0,
// 16'h451c, 16'h4f25, 16'h5790, 16'h5e39,
// 16'h62f4, 16'h65b2, 16'h665f, 16'h64f5,
// 16'h618a, 16'h5c17, 16'h54d1, 16'h4bcd,
// 16'h4142, 16'h3567, 16'h2872, 16'h1aad,
// 16'h0c60, 16'hfdcd, 16'hef51, 16'he11a,
// 16'hd396, 16'hc6e8, 16'hbb70, 16'hb151,
// 16'ha8d2, 16'ha211, 16'h9d3c, 16'h9a65,
// 16'h999e, 16'h9ae8, 16'h9e45, 16'ha392,
// 16'haacb, 16'hb3b3, 16'hbe2e, 16'hc9fc,
// 16'hd6e3, 16'he49d, 16'hf2e8, 16'h0176,
// 16'h0ffa, 16'h1e32, 16'h2bc2, 16'h387c,
// 16'h4405, 16'h4e37, 16'h56cd, 16'h5da3,
// 16'h6292, 16'h6583, 16'h6665, 16'h6534,
// 16'h61f6, 16'h5cb9, 16'h559f, 16'h4cc8,
// 16'h4260, 16'h36a4, 16'h29c7, 16'h1c16,
// 16'h0dd3, 16'hff42, 16'hf0c0, 16'he282,
// 16'hd4e5, 16'hc822, 16'hbc85, 16'hb243,
// 16'ha998, 16'ha2a8, 16'h9da2, 16'h9a95,
// 16'h999a, 16'h9ab1, 16'h9dd5, 16'ha2f7,
// 16'ha9fb, 16'hb2bf, 16'hbd0f, 16'hc8c3,
// 16'hd58a, 16'he33a, 16'hf173, 16'h2002,
// 16'h0e89, 16'h1cca, 16'h2a73, 16'h373f,
// 16'h42ef, 16'h4d42, 16'h5605, 16'h5d0a,
// 16'h622a, 16'h654f, 16'h6668, 16'h6568,
// 16'h6262, 16'h5d53, 16'h566d, 16'h4db9,
// 16'h437f, 16'h37db, 16'h2b1c, 16'h1d7e,
// 16'h0f41, 16'h20bc, 16'hf22f, 16'he3e9,
// 16'hd638, 16'hc95e, 16'hbd9f, 16'hb339,
// 16'haa62, 16'ha343, 16'h9e0e, 16'h9aca,
// 16'h999d, 16'h9a7b, 16'h9d6f, 16'ha25c,
// 16'ha934, 16'hb1ca, 16'hbbf8, 16'hc788,
// 16'hd439, 16'he1d3, 16'hf003, 16'hfe8b,
// 16'h0d19, 16'h1b60, 16'h2920, 16'h3602,
// 16'h41d4, 16'h4c4a, 16'h5539, 16'h5c69,
// 16'h61bf, 16'h6516, 16'h6662, 16'h659c,
// 16'h62c3, 16'h5def, 16'h572f, 16'h4eae,
// 16'h4491, 16'h3916, 16'h2c6e, 16'h1ee0,
// 16'h10b6, 16'h022e, 16'hf3a2, 16'he553,
// 16'hd78b, 16'hca9f, 16'hbeb8, 16'hb437,
// 16'hab2d, 16'ha3e7, 16'h9e7c, 16'h9b05,
// 16'h99a4, 16'h9a4d, 16'h9d0d, 16'ha1c6,
// 16'ha871, 16'hb0da, 16'hbae3, 16'hc653,
// 16'hd2e7, 16'he070, 16'hee92, 16'hfd16,
// 16'h0ba5, 16'h19fa, 16'h27c5, 16'h34c9,
// 16'h40ae, 16'h4b54, 16'h5463, 16'h5bca,
// 16'h614c, 16'h64d8, 16'h6658, 16'h65c7,
// 16'h6325, 16'h5e80, 16'h57f2, 16'h4f99,
// 16'h45a8, 16'h3a47, 16'h2dbf, 16'h2043,
// 16'h1225, 16'h03a6, 16'hf513, 16'he6bc,
// 16'hd8e5, 16'hcbdc, 16'hbfde, 16'hb530,
// 16'hac02, 16'ha48e, 16'h9eed, 16'h9b4b,
// 16'h99ac, 16'h9a26, 16'h9cac, 16'ha13b,
// 16'ha7ad, 16'haff4, 16'hb9ce, 16'hc51f,
// 16'hd19c, 16'hdf0a, 16'hed25, 16'hfba0,
// 16'h0a31, 16'h1890, 16'h266e, 16'h3383,
// 16'h3f91, 16'h4a4f, 16'h5393, 16'h5b1d,
// 16'h60d8, 16'h6493, 16'h664b, 16'h65ee,
// 16'h637d, 16'h5f10, 16'h58ad, 16'h5083,
// 16'h46b8, 16'h3b78, 16'h2f0d, 16'h21a3,
// 16'h1396, 16'h0518, 16'hf68b, 16'he823,
// 16'hda41, 16'hcd1f, 16'hc101, 16'hb633,
// 16'hacd9, 16'ha539, 16'h9f66, 16'h9b90,
// 16'h99bf, 16'h9a01, 16'h9c56, 16'ha0ac,
// 16'ha6f6, 16'haf0a, 16'hb8c4, 16'hc3eb,
// 16'hd053, 16'hdda8, 16'hebb6, 16'hfa2d,
// 16'h08ba, 16'h1729, 16'h250f, 16'h3242,
// 16'h3e67, 16'h494f, 16'h52b7, 16'h5a72,
// 16'h605b, 16'h644a, 16'h6637, 16'h660f,
// 16'h63d4, 16'h5f97, 16'h5966, 16'h5168,
// 16'h47c3, 16'h3ca8, 16'h3056, 16'h2305,
// 16'h1501, 16'h0691, 16'hf7fa, 16'he993,
// 16'hdb9c, 16'hce63, 16'hc22c, 16'hb735,
// 16'hadb7, 16'ha5e6, 16'h9fe7, 16'h9bda,
// 16'h99d5, 16'h99e5, 16'h9bfe, 16'ha02d,
// 16'ha63a, 16'hae2a, 16'hb7b8, 16'hc2c1,
// 16'hcf06, 16'hdc4d, 16'hea45, 16'hf8ba,
// 16'h0746, 16'h15ba, 16'h23b4, 16'h30fa,
// 16'h3d3f, 16'h4847, 16'h51d9, 16'h59c1,
// 16'h5fd8, 16'h63fe, 16'h661e, 16'h662a,
// 16'h6427, 16'h6016, 16'h5a1e, 16'h5246,
// 16'h48cd, 16'h3dd4, 16'h319c, 16'h2465,
// 16'h166d, 16'h0805, 16'hf970, 16'heaff,
// 16'hdcfb, 16'hcfaa, 16'hc358, 16'hb83c,
// 16'hae9a, 16'ha697, 16'ha06d, 16'h9c29,
// 16'h99f2, 16'h99c9, 16'h9bb6, 16'h9fa3,
// 16'ha593, 16'had43, 16'hb6b7, 16'hc194,
// 16'hcdc1, 16'hdaee, 16'he8db, 16'hf742,
// 16'h05d6, 16'h1449, 16'h2257, 16'h2faf,
// 16'h3c13, 16'h473c, 16'h50f7, 16'h590a,
// 16'h5f54, 16'h63a9, 16'h6601, 16'h663e,
// 16'h6473, 16'h6098, 16'h5ac8, 16'h5327,
// 16'h49cd, 16'h3eff, 16'h32e1, 16'h25c0,
// 16'h17db, 16'h0977, 16'hfae6, 16'hec6d,
// 16'hde5a, 16'hd0f5, 16'hc487, 16'hb947,
// 16'haf80, 16'ha74f, 16'ha0f4, 16'h9c80,
// 16'h9a12, 16'h99b8, 16'h9b68, 16'h9f2f,
// 16'ha4dc, 16'hac73, 16'hb5ac, 16'hc073,
// 16'hcc7b, 16'hd993, 16'he770, 16'hf5cf,
// 16'h045e, 16'h12de, 16'h20f4, 16'h2e65,
// 16'h3ae2, 16'h462e, 16'h5010, 16'h5850,
// 16'h5ec8, 16'h6351, 16'h65de, 16'h664e,
// 16'h64bb, 16'h610e, 16'h5b76, 16'h53fc,
// 16'h4ad0, 16'h4022, 16'h3425, 16'h271a,
// 16'h1945, 16'h0aec, 16'hfc59, 16'hedde,
// 16'hdfba, 16'hd244, 16'hc5b6, 16'hba5b,
// 16'hb063, 16'ha812, 16'ha17d, 16'h9cdd,
// 16'h9a39, 16'h99a7, 16'h9b28, 16'h9eb3,
// 16'ha439, 16'hab9a, 16'hb4b0, 16'hbf4e,
// 16'hcb39, 16'hd83a, 16'he608, 16'hf459,
// 16'h02ec, 16'h116c, 16'h1f91, 16'h2d1a,
// 16'h39ab, 16'h4520, 16'h4f22, 16'h5793,
// 16'h5e36, 16'h62f6, 16'h65b2, 16'h665d,
// 16'h64f9, 16'h6185, 16'h5c19, 16'h54d1,
// 16'h4bce, 16'h4142, 16'h3566, 16'h2872,
// 16'h1aad, 16'h0c61, 16'hfdce, 16'hef4c,
// 16'he121, 16'hd38f, 16'hc6ee, 16'hbb6c,
// 16'hb153, 16'ha8d1, 16'ha211, 16'h9d3c,
// 16'h9a65, 16'h999e, 16'h9ae9, 16'h9e42,
// 16'ha396, 16'haac7, 16'hb3b6, 16'hbe2d,
// 16'hc9fb, 16'hd6e4, 16'he49c, 16'hf2ea,
// 16'h0174, 16'h0ffc, 16'h1e2f, 16'h2bc5,
// 16'h3879, 16'h4408, 16'h4e35, 16'h56cd,
// 16'h5da4, 16'h6290, 16'h6586, 16'h6663,
// 16'h6534, 16'h61f6, 16'h5cb8, 16'h55a3,
// 16'h4cc3, 16'h4263, 16'h36a2, 16'h29c9,
// 16'h1c15, 16'h0dd3, 16'hff42, 16'hf0c0,
// 16'he283, 16'hd4e3, 16'hc824, 16'hbc84,
// 16'hb243, 16'ha998, 16'ha2a8, 16'h9da1,
// 16'h9a97, 16'h9998, 16'h9ab2, 16'h9dd4,
// 16'ha2f8, 16'ha9fa, 16'hb2c0, 16'hbd0f,
// 16'hc8c1, 16'hd58e, 16'he335, 16'hf177,
// 16'h2020, 16'h0e89, 16'h1ccb, 16'h2a72,
// 16'h373e, 16'h42f2, 16'h4d3f, 16'h5607,
// 16'h5d08, 16'h622b, 16'h654f, 16'h6668,
// 16'h6568, 16'h6261, 16'h5d55, 16'h566b,
// 16'h4dba, 16'h437f, 16'h37d9, 16'h2b20,
// 16'h1d79, 16'h0f45, 16'h20ba, 16'hf22e,
// 16'he3eb, 16'hd638, 16'hc95c, 16'hbda2,
// 16'hb334, 16'haa67, 16'ha340, 16'h9e10,
// 16'h9ac8, 16'h999f, 16'h9a79, 16'h9d71,
// 16'ha25a, 16'ha935, 16'hb1ca, 16'hbbf8,
// 16'hc788, 16'hd439, 16'he1d3, 16'hf003,
// 16'hfe8b, 16'h0d19, 16'h1b60, 16'h2920,
// 16'h3602, 16'h41d4, 16'h4c4a, 16'h5539,
// 16'h5c6a, 16'h61be, 16'h6516, 16'h6663,
// 16'h659b, 16'h62c4, 16'h5def, 16'h572e,
// 16'h4eae, 16'h4493, 16'h3913, 16'h2c71,
// 16'h1edd, 16'h10b8, 16'h022d, 16'hf3a3,
// 16'he551, 16'hd78e, 16'hca9b, 16'hbebd,
// 16'hb432, 16'hab2f, 16'ha3e9, 16'h9e78,
// 16'h9b09, 16'h99a1, 16'h9a4f, 16'h9d0b,
// 16'ha1c8, 16'ha870, 16'hb0d9, 16'hbae7,
// 16'hc64d, 16'hd2ed, 16'he06c, 16'hee93,
// 16'hfd16, 16'h0ba5, 16'h19fa, 16'h27c6,
// 16'h34c6, 16'h40b1, 16'h4b52, 16'h5464,
// 16'h5bca, 16'h614a, 16'h64da, 16'h6658,
// 16'h65c6, 16'h6326, 16'h5e7f, 16'h57f2,
// 16'h4f9a, 16'h45a6, 16'h3a4a, 16'h2dbb,
// 16'h2047, 16'h1222, 16'h03a8, 16'hf512,
// 16'he6bc, 16'hd8e6, 16'hcbda, 16'hbfe1,
// 16'hb52c, 16'hac07, 16'ha489, 16'h9ef1,
// 16'h9b47, 16'h99af, 16'h9a25, 16'h9cad,
// 16'ha139, 16'ha7af, 16'haff1, 16'hb9d3,
// 16'hc51a, 16'hd1a0, 16'hdf06, 16'hed28,
// 16'hfb9e, 16'h0a34, 16'h188e, 16'h266d,
// 16'h3386, 16'h3f8c, 16'h4a55, 16'h538d,
// 16'h5b23, 16'h60d3, 16'h6496, 16'h6649,
// 16'h65ee, 16'h637f, 16'h5f0f, 16'h58ac,
// 16'h5085, 16'h46b6, 16'h3b7a, 16'h2f0b,
// 16'h21a5, 16'h1394, 16'h051a, 16'hf689,
// 16'he825, 16'hda40, 16'hcd1e, 16'hc104,
// 16'hb62f, 16'hacdd, 16'ha535, 16'h9f69,
// 16'h9b8e, 16'h99c1, 16'h99ff, 16'h9c57,
// 16'ha0ac, 16'ha6f7, 16'haf08, 16'hb8c4,
// 16'hc3ee, 16'hd050, 16'hdda9, 16'hebb7,
// 16'hfa29, 16'h08c1, 16'h1722, 16'h2513,
// 16'h323f, 16'h3e6a, 16'h494d, 16'h52b9,
// 16'h5a70, 16'h605b, 16'h644b, 16'h6637,
// 16'h660e, 16'h63d6, 16'h5f94, 16'h596a,
// 16'h5164, 16'h47c6, 16'h3ca7, 16'h3055,
// 16'h2308, 16'h14fe, 16'h0692, 16'hf7fb,
// 16'he992, 16'hdb9c, 16'hce64, 16'hc22a,
// 16'hb736, 16'hadb7, 16'ha5e6, 16'h9fe6,
// 16'h9bdb, 16'h99d5, 16'h99e3, 16'h9c02,
// 16'ha027, 16'ha640, 16'hae26, 16'hb7ba,
// 16'hc2c0, 16'hcf07, 16'hdc4b, 16'hea48,
// 16'hf8b6, 16'h074b, 16'h15b6, 16'h23b8,
// 16'h30f6, 16'h3d41, 16'h4847, 16'h51d9,
// 16'h59c1, 16'h5fd8, 16'h63fd, 16'h661f,
// 16'h6629, 16'h6427, 16'h6018, 16'h5a1b,
// 16'h5247, 16'h48cd, 16'h3dd2, 16'h31a0,
// 16'h2461, 16'h1670, 16'h0802, 16'hf973,
// 16'heafc, 16'hdcfe, 16'hcfa7, 16'hc35a,
// 16'hb83c, 16'hae99, 16'ha699, 16'ha06b,
// 16'h9c29, 16'h99f3, 16'h99ca, 16'h9bb3,
// 16'h9fa7, 16'ha58e, 16'had47, 16'hb6b5,
// 16'hc195, 16'hcdc1, 16'hdaed, 16'he8dd,
// 16'hf740, 16'h05d7, 16'h1449, 16'h2257,
// 16'h2faf, 16'h3c13, 16'h473c, 16'h50f8,
// 16'h5908, 16'h5f55, 16'h63a9, 16'h6620,
// 16'h6640, 16'h6471, 16'h6098, 16'h5aca,
// 16'h5324, 16'h49d0, 16'h3efd, 16'h32e1,
// 16'h25c2, 16'h17d8, 16'h097a, 16'hfae4,
// 16'hec6e, 16'hde59, 16'hd0f6, 16'hc486,
// 16'hb949, 16'haf7d, 16'ha752, 16'ha0f2,
// 16'h9c81, 16'h9a13, 16'h99b5, 16'h9b6c,
// 16'h9f2b, 16'ha4df, 16'hac71, 16'hb5ae,
// 16'hc071, 16'hcc7d, 16'hd990, 16'he774,
// 16'hf5cb, 16'h0463, 16'h12d8, 16'h20f9,
// 16'h2e62, 16'h3ae3, 16'h4630, 16'h500c,
// 16'h5854, 16'h5ec4, 16'h6356, 16'h65d8,
// 16'h6654, 16'h64b6, 16'h6112, 16'h5b74,
// 16'h53fc, 16'h4ad1, 16'h4022, 16'h3423,
// 16'h271e, 16'h1941, 16'h0aed, 16'hfc5b,
// 16'heddb, 16'hdfbd, 16'hd242, 16'hc5b6,
// 16'hba5b, 16'hb065, 16'ha80f, 16'ha181,
// 16'h9cd9, 16'h9a3c, 16'h99a5, 16'h9b29,
// 16'h9eb4, 16'ha437, 16'hab9b, 16'hb4b0,
// 16'hbf4c, 16'hcb3d, 16'hd836, 16'he60a,
// 16'hf458, 16'h02ec, 16'h116c, 16'h1f92,
// 16'h2d17, 16'h39af, 16'h451c, 16'h4f26,
// 16'h578e, 16'h5e3b, 16'h62f3, 16'h65b2,
// 16'h6660, 16'h64f4, 16'h618a, 16'h5c17,
// 16'h54d1, 16'h4bcd, 16'h4144, 16'h3563,
// 16'h2875, 16'h1aac, 16'h0c60, 16'hfdcf,
// 16'hef4c, 16'he11f, 16'hd393, 16'hc6eb,
// 16'hbb6d, 16'hb153, 16'ha8d0, 16'ha213,
// 16'h9d3b, 16'h9a65, 16'h999d, 16'h9aeb,
// 16'h9e41, 16'ha396, 16'haac8, 16'hb3b4,
// 16'hbe2e, 16'hc9fd, 16'hd6e1, 16'he4a0,
// 16'hf2e6, 16'h0176, 16'h0ffb, 16'h1e30,
// 16'h2bc5, 16'h3879, 16'h4408, 16'h4e35,
// 16'h56cd, 16'h5da3, 16'h6293, 16'h6581,
// 16'h666a, 16'h652d, 16'h61fb, 16'h5cb6,
// 16'h55a2, 16'h4cc6, 16'h4261, 16'h36a3,
// 16'h29c7, 16'h1c17, 16'h0dd1, 16'hff45,
// 16'hf0be, 16'he283, 16'hd4e3, 16'hc824,
// 16'hbc84, 16'hb244, 16'ha997, 16'ha2a8,
// 16'h9da3, 16'h9a93, 16'h999d, 16'h9aae,
// 16'h9dd6, 16'ha2f7, 16'ha9fb, 16'hb2be,
// 16'hbd12, 16'hc8be, 16'hd58f, 16'he336,
// 16'hf176, 16'h2001, 16'h0e88, 16'h1ccc,
// 16'h2a70, 16'h3742, 16'h42ed, 16'h4d44,
// 16'h5603, 16'h5d0b, 16'h6229, 16'h6550,
// 16'h6666, 16'h656b, 16'h625e, 16'h5d59,
// 16'h5666, 16'h4dc0, 16'h4378, 16'h37e0,
// 16'h2b1b, 16'h1d7c, 16'h0f44, 16'h20ba,
// 16'hf22f, 16'he3eb, 16'hd636, 16'hc95f,
// 16'hbd9e, 16'hb33a, 16'haa60, 16'ha347,
// 16'h9e09, 16'h9ace, 16'h999b, 16'h9a7c,
// 16'h9d6f, 16'ha25b, 16'ha935, 16'hb1ca,
// 16'hbbf8, 16'hc789, 16'hd437, 16'he1d5,
// 16'hf001, 16'hfe8d, 16'h0d17, 16'h1b62,
// 16'h291e, 16'h3604, 16'h41d3, 16'h4c49,
// 16'h553a, 16'h5c69, 16'h61c1, 16'h6513,
// 16'h6665, 16'h6598, 16'h62c8, 16'h5dec,
// 16'h572f, 16'h4eaf, 16'h4490, 16'h3917,
// 16'h2c6e, 16'h1edf, 16'h10b6, 16'h022e,
// 16'hf3a3, 16'he551, 16'hd78f, 16'hca99,
// 16'hbebe, 16'hb432, 16'hab30, 16'ha3e6,
// 16'h9e7c, 16'h9b05, 16'h99a5, 16'h9a4c,
// 16'h9d0c, 16'ha1c8, 16'ha870, 16'hb0da,
// 16'hbae5, 16'hc650, 16'hd2e9, 16'he06f,
// 16'hee92, 16'hfd17, 16'h0ba4, 16'h19fb,
// 16'h27c5, 16'h34c6, 16'h40b3, 16'h4b4f,
// 16'h5468, 16'h5bc6, 16'h614d, 16'h64d8,
// 16'h6658, 16'h65c9, 16'h6322, 16'h5e82,
// 16'h57f1, 16'h4f99, 16'h45a8, 16'h3a48,
// 16'h2dbd, 16'h2046, 16'h1222, 16'h03a8,
// 16'hf512, 16'he6bb, 16'hd8e7, 16'hcbda,
// 16'hbfe0, 16'hb52f, 16'hac02, 16'ha48d,
// 16'h9eef, 16'h9b48, 16'h99af, 16'h9a25,
// 16'h9cad, 16'ha139, 16'ha7af, 16'haff1,
// 16'hb9d2, 16'hc51d, 16'hd19c, 16'hdf0b,
// 16'hed24, 16'hfba0, 16'h0a32, 16'h188f,
// 16'h266f, 16'h3383, 16'h3f8f, 16'h4a51,
// 16'h5391, 16'h5b20, 16'h60d5, 16'h6495,
// 16'h6649, 16'h65ef, 16'h637e, 16'h5f0e,
// 16'h58af, 16'h5082, 16'h46b8, 16'h3b79,
// 16'h2f0b, 16'h21a6, 16'h1393, 16'h051b,
// 16'hf687, 16'he827, 16'hda3f, 16'hcd1f,
// 16'hc102, 16'hb630, 16'hacdd, 16'ha535,
// 16'h9f69, 16'h9b8f, 16'h99be, 16'h9a03,
// 16'h9c54, 16'ha0ae, 16'ha6f5, 16'haf0a,
// 16'hb8c3, 16'hc3ee, 16'hd050, 16'hdda9,
// 16'hebb7, 16'hfa29, 16'h08c2, 16'h171f,
// 16'h2517, 16'h323c, 16'h3e6c, 16'h494d,
// 16'h52b5, 16'h5a75, 16'h6058, 16'h644d,
// 16'h6636, 16'h660e, 16'h63d5, 16'h5f97,
// 16'h5965, 16'h516b, 16'h47be, 16'h3caf,
// 16'h304e, 16'h230c, 16'h14fd, 16'h0692,
// 16'hf7fc, 16'he990, 16'hdb9e, 16'hce62,
// 16'hc22c, 16'hb736, 16'hadb6, 16'ha5e6,
// 16'h9fe7, 16'h9bd9, 16'h99d7, 16'h99e2,
// 16'h9c02, 16'ha028, 16'ha63f, 16'hae26,
// 16'hb7ba, 16'hc2c0, 16'hcf09, 16'hdc48,
// 16'hea4b, 16'hf8b3, 16'h074d, 16'h15b5,
// 16'h23b9, 16'h30f4, 16'h3d44, 16'h4843,
// 16'h51db, 16'h59c1, 16'h5fd8, 16'h63fe,
// 16'h661d, 16'h662b, 16'h6424, 16'h601c,
// 16'h5a18, 16'h524a, 16'h48cb, 16'h3dd2,
// 16'h31a1, 16'h245f, 16'h1673, 16'h0820,
// 16'hf973, 16'heafd, 16'hdcfc, 16'hcfa9,
// 16'hc359, 16'hb83c, 16'hae99, 16'ha699,
// 16'ha06a, 16'h9c2b, 16'h99f1, 16'h99cb,
// 16'h9bb3, 16'h9fa7, 16'ha58e, 16'had48,
// 16'hb6b3, 16'hc196, 16'hcdc2, 16'hdaec,
// 16'he8dd, 16'hf741, 16'h05d5, 16'h144b,
// 16'h2255, 16'h2fb2, 16'h3c10, 16'h473e,
// 16'h50f6, 16'h590a, 16'h5f54, 16'h63aa,
// 16'h65fe, 16'h6643, 16'h646f, 16'h6098,
// 16'h5acb, 16'h5323, 16'h49d1, 16'h3efc,
// 16'h32e2, 16'h25c1, 16'h17da, 16'h0977,
// 16'hfae6, 16'hec6d, 16'hde5a, 16'hd0f6,
// 16'hc484, 16'hb94c, 16'haf7a, 16'ha755,
// 16'ha0ef, 16'h9c84, 16'h9a10, 16'h99b7,
// 16'h9b6b, 16'h9f2a, 16'ha4e3, 16'hac6c,
// 16'hb5b1, 16'hc070, 16'hcc7c, 16'hd993,
// 16'he770, 16'hf5ce, 16'h0460, 16'h12dc,
// 16'h20f5, 16'h2e65, 16'h3ae1, 16'h462f,
// 16'h5010, 16'h584e, 16'h5ecb, 16'h634f,
// 16'h65de, 16'h6650, 16'h64b8, 16'h6110,
// 16'h5b77, 16'h53f9, 16'h4ad4, 16'h401e,
// 16'h3428, 16'h2718, 16'h1948, 16'h0ae7,
// 16'hfc5f, 16'hedd9, 16'hdfbd, 16'hd243,
// 16'hc5b5, 16'hba5c, 16'hb065, 16'ha80e,
// 16'ha182, 16'h9cd8, 16'h9a3d, 16'h99a4,
// 16'h9b2b, 16'h9eb1, 16'ha43b, 16'hab97,
// 16'hb4b2, 16'hbf4d, 16'hcb3b, 16'hd839,
// 16'he606, 16'hf45c, 16'h02e9, 16'h116e,
// 16'h1f92, 16'h2d16, 16'h39af, 16'h451c,
// 16'h4f26, 16'h578f, 16'h5e3a, 16'h62f3,
// 16'h65b2, 16'h6660, 16'h64f4, 16'h618a,
// 16'h5c17, 16'h54d1, 16'h4bce, 16'h4142,
// 16'h3566, 16'h2871, 16'h1ab0, 16'h0c5c,
// 16'hfdd3, 16'hef4a, 16'he120, 16'hd390,
// 16'hc6ef, 16'hbb69, 16'hb157, 16'ha8cd,
// 16'ha215, 16'h9d39, 16'h9a67, 16'h999c,
// 16'h9aeb, 16'h9e42, 16'ha393, 16'haacc,
// 16'hb3b1, 16'hbe30, 16'hc9fc, 16'hd6e0,
// 16'he4a1, 16'hf2e5, 16'h0178, 16'h0ff9,
// 16'h1e32, 16'h2bc2, 16'h387c, 16'h4405,
// 16'h4e37, 16'h56cd, 16'h5da3, 16'h6291,
// 16'h6585, 16'h6663, 16'h6536, 16'h61f3,
// 16'h5cbc, 16'h559e, 16'h4cc7, 16'h4262,
// 16'h36a1, 16'h29cb, 16'h1c13, 16'h0dd3,
// 16'hff45, 16'hf0bd, 16'he284, 16'hd4e3,
// 16'hc824, 16'hbc84, 16'hb245, 16'ha994,
// 16'ha2ac, 16'h9d9e, 16'h9a99, 16'h9998,
// 16'h9ab1, 16'h9dd6, 16'ha2f4, 16'ha9ff,
// 16'hb2bb, 16'hbd13, 16'hc8bf, 16'hd58e,
// 16'he336, 16'hf177, 16'hfffe, 16'h0e8c,
// 16'h1cc8, 16'h2a74, 16'h373f, 16'h42ef,
// 16'h4d41, 16'h5607, 16'h5d06, 16'h622f,
// 16'h654c, 16'h6668, 16'h6569, 16'h6260,
// 16'h5d57, 16'h5668, 16'h4dbf, 16'h4377,
// 16'h37e3, 16'h2b17, 16'h1d80, 16'h0f40,
// 16'h20bd, 16'hf22d, 16'he3ec, 16'hd636,
// 16'hc95f, 16'hbd9e, 16'hb339, 16'haa62,
// 16'ha344, 16'h9e0d, 16'h9aca, 16'h999d,
// 16'h9a7c, 16'h9d6e, 16'ha25d, 16'ha933,
// 16'hb1c9, 16'hbbfb, 16'hc785, 16'hd43d,
// 16'he1cf, 16'hf005, 16'hfe8a, 16'h0d19,
// 16'h1b62, 16'h291e, 16'h3603, 16'h41d4,
// 16'h4c49, 16'h5539, 16'h5c6b, 16'h61bd,
// 16'h6517, 16'h6662, 16'h659b, 16'h62c4,
// 16'h5df0, 16'h572c, 16'h4eb0, 16'h4491,
// 16'h3916, 16'h2c6d, 16'h1ee2, 16'h10b3,
// 16'h0231, 16'hf3a0, 16'he554, 16'hd78b,
// 16'hca9e, 16'hbeba, 16'hb435, 16'hab2e,
// 16'ha3e8, 16'h9e79, 16'h9b08, 16'h99a2,
// 16'h9a4f, 16'h9d0a, 16'ha1c9, 16'ha86f,
// 16'hb0db, 16'hbae4, 16'hc650, 16'hd2eb,
// 16'he06c, 16'hee95, 16'hfd14, 16'h0ba7,
// 16'h19f8, 16'h27c8, 16'h34c4, 16'h40b3,
// 16'h4b50, 16'h5466, 16'h5bc9, 16'h614b,
// 16'h64d8, 16'h6659, 16'h65c6, 16'h6326,
// 16'h5e7f, 16'h57f3, 16'h4f98, 16'h45a8,
// 16'h3a47, 16'h2dc0, 16'h2042, 16'h1227,
// 16'h03a2, 16'hf516, 16'he6bb, 16'hd8e6,
// 16'hcbdb, 16'hbfde, 16'hb530, 16'hac03,
// 16'ha48c, 16'h9eef, 16'h9b49, 16'h99ad,
// 16'h9a27, 16'h9cab, 16'ha13b, 16'ha7ae,
// 16'haff1, 16'hb9d2, 16'hc51d, 16'hd19d,
// 16'hdf09, 16'hed26, 16'hfb9e, 16'h0a34,
// 16'h188e, 16'h266e, 16'h3384, 16'h3f8f,
// 16'h4a51, 16'h5391, 16'h5b1f, 16'h60d7,
// 16'h6492, 16'h664d, 16'h65eb, 16'h6382,
// 16'h5f0a, 16'h58b2, 16'h5080, 16'h46b9,
// 16'h3b79, 16'h2f0a, 16'h21a7, 16'h1391,
// 16'h051e, 16'hf684, 16'he829, 16'hda3e,
// 16'hcd1e, 16'hc104, 16'hb62f, 16'hacde,
// 16'ha533, 16'h9f6b, 16'h9b8c, 16'h99c2,
// 16'h99ff, 16'h9c57, 16'ha0ac, 16'ha6f7,
// 16'haf07, 16'hb8c6, 16'hc3eb, 16'hd053,
// 16'hdda8, 16'hebb7, 16'hfa29, 16'h08c0,
// 16'h1723, 16'h2513, 16'h3240, 16'h3e68,
// 16'h494e, 16'h52b9, 16'h5a6f, 16'h605e,
// 16'h6447, 16'h663a, 16'h660d, 16'h63d5,
// 16'h5f97, 16'h5965, 16'h516a, 16'h47c0,
// 16'h3cab, 16'h3054, 16'h2306, 16'h1501,
// 16'h0690, 16'hf7fc, 16'he991, 16'hdb9d,
// 16'hce63, 16'hc22b, 16'hb736, 16'hadb7,
// 16'ha5e5, 16'h9fe9, 16'h9bd7, 16'h99d8,
// 16'h99e2, 16'h9c01, 16'ha02b, 16'ha63b,
// 16'hae2a, 16'hb7b7, 16'hc2c2, 16'hcf07,
// 16'hdc4a, 16'hea49, 16'hf8b6, 16'h0749,
// 16'h15ba, 16'h23b1, 16'h30fe, 16'h3d3b,
// 16'h484b, 16'h51d6, 16'h59c2, 16'h5fd8,
// 16'h63fe, 16'h661f, 16'h6628, 16'h6428,
// 16'h6016, 16'h5a1f, 16'h5245, 16'h48ce,
// 16'h3dd1, 16'h319f, 16'h2463, 16'h166e,
// 16'h0806, 16'hf96d, 16'heb02, 16'hdcf7,
// 16'hcfae, 16'hc355, 16'hb83f, 16'hae96,
// 16'ha69c, 16'ha068, 16'h9c2c, 16'h99f1,
// 16'h99c9, 16'h9bb5, 16'h9fa7, 16'ha58c,
// 16'had4a, 16'hb6b1, 16'hc198, 16'hcdc0,
// 16'hdaed, 16'he8de, 16'hf73e, 16'h05da,
// 16'h1445, 16'h225b, 16'h2fad, 16'h3c13,
// 16'h473e, 16'h50f3, 16'h590e, 16'h5f51,
// 16'h63ac, 16'h65fe, 16'h6641, 16'h6470,
// 16'h609a, 16'h5ac7, 16'h5327, 16'h49cf,
// 16'h3efc, 16'h32e3, 16'h25bf, 16'h17db,
// 16'h0977, 16'hfae8, 16'hec69, 16'hde5e,
// 16'hd0f2, 16'hc488, 16'hb949, 16'haf7d,
// 16'ha751, 16'ha0f4, 16'h9c7e, 16'h9a16,
// 16'h99b3, 16'h9b6c, 16'h9f2c, 16'ha4df,
// 16'hac70, 16'hb5af, 16'hc06f, 16'hcc7f,
// 16'hd990, 16'he773, 16'hf5ca, 16'h0464,
// 16'h12da, 16'h20f6, 16'h2e64, 16'h3ae1,
// 16'h4630, 16'h500f, 16'h5851, 16'h5ec6,
// 16'h6354, 16'h65d9, 16'h6654, 16'h64b7,
// 16'h6110, 16'h5b75, 16'h53fd, 16'h4ace,
// 16'h4026, 16'h3421, 16'h271c, 16'h1945,
// 16'h0aea, 16'hfc5d, 16'hedda, 16'hdfbd,
// 16'hd242, 16'hc5b6, 16'hba5c, 16'hb063,
// 16'ha812, 16'ha17d, 16'h9cdd, 16'h9a39,
// 16'h99a6, 16'h9b2a, 16'h9eb2, 16'ha43a,
// 16'hab98, 16'hb4b0, 16'hbf4f, 16'hcb39,
// 16'hd83b, 16'he605, 16'hf45b, 16'h02ec,
// 16'h116b, 16'h1f93, 16'h2d17, 16'h39ad,
// 16'h4520, 16'h4f22, 16'h5792, 16'h5e37,
// 16'h62f6, 16'h65b1, 16'h665e, 16'h64f9,
// 16'h6184, 16'h5c1c, 16'h54ce, 16'h4bce,
// 16'h4144, 16'h3563, 16'h2875, 16'h1aab,
// 16'h0c62, 16'hfdcd, 16'hef4e, 16'he11e,
// 16'hd392, 16'hc6eb, 16'hbb6f, 16'hb151,
// 16'ha8d2, 16'ha210, 16'h9d3e, 16'h9a62,
// 16'h99a2, 16'h9ae5, 16'h9e46, 16'ha393,
// 16'haac9, 16'hb3b5, 16'hbe2d, 16'hc9fd,
// 16'hd6e1, 16'he4a0, 16'hf2e5, 16'h0178,
// 16'h0ffa, 16'h1e30, 16'h2bc5, 16'h3879,
// 16'h4407, 16'h4e37, 16'h56cb, 16'h5da6,
// 16'h628f, 16'h6586, 16'h6662, 16'h6536,
// 16'h61f4, 16'h5cba, 16'h55a1, 16'h4cc4,
// 16'h4263, 16'h36a2, 16'h29c7, 16'h1c18,
// 16'h0dd0, 16'hff45, 16'hf0bf, 16'he281,
// 16'hd4e7, 16'hc820, 16'hbc86, 16'hb244,
// 16'ha996, 16'ha2ab, 16'h9d9e, 16'h9a98,
// 16'h9999, 16'h9ab1, 16'h9dd5, 16'ha2f7,
// 16'ha9fa, 16'hb2c0, 16'hbd0f, 16'hc8c1,
// 16'hd58e, 16'he335, 16'hf178, 16'hfffe,
// 16'h0e8b, 16'h1cc9, 16'h2a73, 16'h373f,
// 16'h42f1, 16'h4d3f, 16'h5608, 16'h5d05,
// 16'h6230, 16'h654a, 16'h666b, 16'h6567,
// 16'h625f, 16'h5d5a, 16'h5665, 16'h4dc0,
// 16'h437a, 16'h37dd, 16'h2b1c, 16'h1d7d,
// 16'h0f42, 16'h20bc, 16'hf22e, 16'he3ea,
// 16'hd638, 16'hc95d, 16'hbda0, 16'hb338,
// 16'haa61, 16'ha347, 16'h9e09, 16'h9ace,
// 16'h999a, 16'h9a7d, 16'h9d6f, 16'ha25b,
// 16'ha934, 16'hb1cb, 16'hbbf7, 16'hc789,
// 16'hd439, 16'he1d1, 16'hf006, 16'hfe89,
// 16'h0d19, 16'h1b62, 16'h291d, 16'h3605,
// 16'h41d2, 16'h4c4b, 16'h5538, 16'h5c6a,
// 16'h61bf, 16'h6516, 16'h6662, 16'h659c,
// 16'h62c2, 16'h5df1, 16'h572d, 16'h4eaf,
// 16'h4491, 16'h3916, 16'h2c6d, 16'h1ee2,
// 16'h10b3, 16'h0230, 16'hf3a2, 16'he551,
// 16'hd78f, 16'hca99, 16'hbec0, 16'hb42f,
// 16'hab33, 16'ha3e4, 16'h9e7c, 16'h9b06,
// 16'h99a5, 16'h9a4b, 16'h9d0e, 16'ha1c6,
// 16'ha86f, 16'hb0de, 16'hbae1, 16'hc651,
// 16'hd2ec, 16'he06a, 16'hee97, 16'hfd14,
// 16'h0ba5, 16'h19fa, 16'h27c6, 16'h34c5,
// 16'h40b5, 16'h4b4d, 16'h5469, 16'h5bc5,
// 16'h614e, 16'h64d7, 16'h665a, 16'h65c6,
// 16'h6326, 16'h5e7e, 16'h57f4, 16'h4f97,
// 16'h45a9, 16'h3a48, 16'h2dbe, 16'h2043,
// 16'h1226, 16'h03a3, 16'hf517, 16'he6ba,
// 16'hd8e6, 16'hcbdb, 16'hbfdf, 16'hb52f,
// 16'hac04, 16'ha48c, 16'h9eee, 16'h9b4b,
// 16'h99ab, 16'h9a27, 16'h9cad, 16'ha138,
// 16'ha7b2, 16'hafed, 16'hb9d4, 16'hc51c,
// 16'hd19d, 16'hdf0a, 16'hed25, 16'hfb9e,
// 16'h0a34, 16'h188e, 16'h266d, 16'h3386,
// 16'h3f8d, 16'h4a53, 16'h538e, 16'h5b23,
// 16'h60d1, 16'h6499, 16'h6647, 16'h65ef,
// 16'h637f, 16'h5f0d, 16'h58b0, 16'h5081,
// 16'h46b8, 16'h3b79, 16'h2f0c, 16'h21a5,
// 16'h1394, 16'h051a, 16'hf687, 16'he827,
// 16'hda40, 16'hcd1d, 16'hc105, 16'hb62e,
// 16'hacdd, 16'ha535, 16'h9f6a, 16'h9b8d,
// 16'h99c1, 16'h99ff, 16'h9c57, 16'ha0ad,
// 16'ha6f4, 16'haf0b, 16'hb8c3, 16'hc3ee,
// 16'hd04f, 16'hddab, 16'hebb4, 16'hfa2e,
// 16'h08bc, 16'h1725, 16'h2512, 16'h3240,
// 16'h3e69, 16'h494f, 16'h52b5, 16'h5a74,
// 16'h6058, 16'h644e, 16'h6634, 16'h6611,
// 16'h63d2, 16'h5f99, 16'h5965, 16'h5169,
// 16'h47c2, 16'h3ca9, 16'h3055, 16'h2307,
// 16'h14ff, 16'h0692, 16'hf7fa, 16'he993,
// 16'hdb9c, 16'hce63, 16'hc22b, 16'hb736,
// 16'hadb6, 16'ha5e7, 16'h9fe7, 16'h9bd8,
// 16'h99d8, 16'h99e1, 16'h9c03, 16'ha028,
// 16'ha63d, 16'hae29, 16'hb7b8, 16'hc2c1,
// 16'hcf07, 16'hdc4a, 16'hea4a, 16'hf8b4,
// 16'h074c, 16'h15b6, 16'h23b6, 16'h30fa,
// 16'h3d3d, 16'h484a, 16'h51d6, 16'h59c3,
// 16'h5fd8, 16'h63fd, 16'h6620, 16'h6626,
// 16'h642b, 16'h6014, 16'h5a1f, 16'h5245,
// 16'h48ce, 16'h3dd2, 16'h319f, 16'h2462,
// 16'h166f, 16'h0804, 16'hf971, 16'heaff,
// 16'hdcf9, 16'hcfac, 16'hc357, 16'hb83d,
// 16'hae9a, 16'ha697, 16'ha06c, 16'h9c29,
// 16'h99f3, 16'h99c8, 16'h9bb7, 16'h9fa3,
// 16'ha591, 16'had46, 16'hb6b4, 16'hc196,
// 16'hcdc1, 16'hdaed, 16'he8dd, 16'hf741,
// 16'h05d5, 16'h144b, 16'h2255, 16'h2fb2,
// 16'h3c10, 16'h473f, 16'h50f4, 16'h590c,
// 16'h5f53, 16'h63aa, 16'h65ff, 16'h6641,
// 16'h6470, 16'h609a, 16'h5ac7, 16'h5327,
// 16'h49ce, 16'h3efe, 16'h32e0, 16'h25c4,
// 16'h17d5, 16'h097e, 16'hfae0, 16'hec70,
// 16'hde59, 16'hd0f6, 16'hc486, 16'hb948,
// 16'haf7f, 16'ha750, 16'ha0f4, 16'h9c80,
// 16'h9a12, 16'h99b7, 16'h9b6a, 16'h9f2c,
// 16'ha4e0, 16'hac6f, 16'hb5b0, 16'hc06f,
// 16'hcc7d, 16'hd992, 16'he771, 16'hf5ce,
// 16'h0460, 16'h12db, 16'h20f6, 16'h2e64,
// 16'h3ae2, 16'h462f, 16'h500f, 16'h5851,
// 16'h5ec7, 16'h6352, 16'h65dc, 16'h6651,
// 16'h64b8, 16'h6110, 16'h5b76, 16'h53fa,
// 16'h4ad4, 16'h401d, 16'h3429, 16'h2718,
// 16'h1946, 16'h0aeb, 16'hfc5a, 16'heddd,
// 16'hdfbc, 16'hd241, 16'hc5b9, 16'hba58,
// 16'hb066, 16'ha80f, 16'ha180, 16'h9cdb,
// 16'h9a39, 16'h99a8, 16'h9b26, 16'h9eb7,
// 16'ha435, 16'hab9c, 16'hb4ae, 16'hbf50,
// 16'hcb39, 16'hd83a, 16'he606, 16'hf45b,
// 16'h02eb, 16'h116d, 16'h1f91, 16'h2d17,
// 16'h39af, 16'h451d, 16'h4f26, 16'h578e,
// 16'h5e3a, 16'h62f3, 16'h65b4, 16'h665d,
// 16'h64f8, 16'h6186, 16'h5c18, 16'h54d4,
// 16'h4bc9, 16'h4147, 16'h3561, 16'h2875,
// 16'h1aae, 16'h0c5e, 16'hfdd1, 16'hef4b,
// 16'he11e, 16'hd394, 16'hc6ea, 16'hbb6f,
// 16'hb151, 16'ha8d2, 16'ha210, 16'h9d3e,
// 16'h9a63, 16'h999f, 16'h9ae9, 16'h9e42,
// 16'ha395, 16'haac9, 16'hb3b4, 16'hbe2e,
// 16'hc9fc, 16'hd6e2, 16'he49f, 16'hf2e6,
// 16'h0177, 16'h0ffb, 16'h1e2f, 16'h2bc6,
// 16'h3877, 16'h440b, 16'h4e32, 16'h56cf,
// 16'h5da2, 16'h6293, 16'h6583, 16'h6665,
// 16'h6533, 16'h61f6, 16'h5cba, 16'h559f,
// 16'h4cc7, 16'h4261, 16'h36a2, 16'h29ca,
// 16'h1c14, 16'h0dd2, 16'hff46, 16'hf0bb,
// 16'he287, 16'hd4e1, 16'hc824, 16'hbc85,
// 16'hb243, 16'ha997, 16'ha2a9, 16'h9da1,
// 16'h9a96, 16'h999b, 16'h9aaf, 16'h9dd6,
// 16'ha2f6, 16'ha9fc, 16'hb2be, 16'hbd12,
// 16'hc8bf, 16'hd58e, 16'he336, 16'hf176,
// 16'h2020, 16'h0e8b, 16'h1cc9, 16'h2a72,
// 16'h3740, 16'h42ef, 16'h4d42, 16'h5605,
// 16'h5d09, 16'h622b, 16'h654f, 16'h6668,
// 16'h6567, 16'h6262, 16'h5d55, 16'h566a,
// 16'h4dbd, 16'h437b, 16'h37dd, 16'h2b1d,
// 16'h1d7b, 16'h0f44, 16'h20ba, 16'hf231,
// 16'he3e7, 16'hd63a, 16'hc95c, 16'hbda0,
// 16'hb339, 16'haa61, 16'ha344, 16'h9e0d,
// 16'h9acb, 16'h999c, 16'h9a7c, 16'h9d6e,
// 16'ha25c, 16'ha935, 16'hb1c9, 16'hbbf9,
// 16'hc787, 16'hd43a, 16'he1d1, 16'hf006,
// 16'hfe88, 16'h0d1b, 16'h1b60, 16'h291f,
// 16'h3603, 16'h41d3, 16'h4c4b, 16'h5538,
// 16'h5c6b, 16'h61bd, 16'h6518, 16'h6660,
// 16'h659e, 16'h62c2, 16'h5def, 16'h572f,
// 16'h4ead, 16'h4495, 16'h3911, 16'h2c71,
// 16'h1edf, 16'h10b5, 16'h0231, 16'hf39f,
// 16'he553, 16'hd78e, 16'hca9a, 16'hbebf,
// 16'hb430, 16'hab31, 16'ha3e7, 16'h9e79,
// 16'h9b08, 16'h99a4, 16'h9a4b, 16'h9d0f,
// 16'ha1c5, 16'ha870, 16'hb0dc, 16'hbae3,
// 16'hc651, 16'hd2ea, 16'he06d, 16'hee94,
// 16'hfd15, 16'h0ba6, 16'h19f9, 16'h27c6,
// 16'h34c7, 16'h40b1, 16'h4b50, 16'h5468,
// 16'h5bc6, 16'h614d, 16'h64d7, 16'h665a,
// 16'h65c6, 16'h6326, 16'h5e7f, 16'h57f1,
// 16'h4f9b, 16'h45a6, 16'h3a49, 16'h2dbe,
// 16'h2044, 16'h1224, 16'h03a6, 16'hf514,
// 16'he6bb, 16'hd8e6, 16'hcbdb, 16'hbfde,
// 16'hb531, 16'hac01, 16'ha48e, 16'h9eed,
// 16'h9b4a, 16'h99ad, 16'h9a26, 16'h9cad,
// 16'ha139, 16'ha7af, 16'haff1, 16'hb9d1,
// 16'hc51f, 16'hd19a, 16'hdf0d, 16'hed22,
// 16'hfba2, 16'h0a30, 16'h1891, 16'h266c,
// 16'h3386, 16'h3f8d, 16'h4a53, 16'h5390,
// 16'h5b1f, 16'h60d7, 16'h6491, 16'h6650,
// 16'h65e7, 16'h6386, 16'h5f07, 16'h58b4,
// 16'h507f, 16'h46b9, 16'h3b79, 16'h2f0b,
// 16'h21a6, 16'h1393, 16'h051b, 16'hf687,
// 16'he827, 16'hda3f, 16'hcd1e, 16'hc104,
// 16'hb62f, 16'hacdd, 16'ha535, 16'h9f69,
// 16'h9b8e, 16'h99c1, 16'h99ff, 16'h9c58,
// 16'ha0ab, 16'ha6f7, 16'haf09, 16'hb8c4,
// 16'hc3ed, 16'hd050, 16'hddaa, 16'hebb7,
// 16'hfa29, 16'h08c0, 16'h1722, 16'h2514,
// 16'h3240, 16'h3e67, 16'h4950, 16'h52b6,
// 16'h5a74, 16'h6057, 16'h644f, 16'h6632,
// 16'h6613, 16'h63d3, 16'h5f96, 16'h5967,
// 16'h5168, 16'h47c2, 16'h3cab, 16'h3052,
// 16'h2309, 16'h14fe, 16'h0692, 16'hf7fb,
// 16'he991, 16'hdb9f, 16'hce5f, 16'hc22f,
// 16'hb733, 16'hadb8, 16'ha5e7, 16'h9fe4,
// 16'h9bdc, 16'h99d6, 16'h99e1, 16'h9c04,
// 16'ha027, 16'ha63e, 16'hae29, 16'hb7b6,
// 16'hc2c4, 16'hcf04, 16'hdc4d, 16'hea47,
// 16'hf8b7, 16'h0749, 16'h15b9, 16'h23b3,
// 16'h30fb, 16'h3d3f, 16'h4847, 16'h51d9,
// 16'h59c0, 16'h5fda, 16'h63fd, 16'h661e,
// 16'h662a, 16'h6425, 16'h601b, 16'h5a19,
// 16'h5249, 16'h48cb, 16'h3dd5, 16'h319c,
// 16'h2465, 16'h166c, 16'h0807, 16'hf96d,
// 16'heb02, 16'hdcf9, 16'hcfaa, 16'hc359,
// 16'hb83b, 16'hae9b, 16'ha697, 16'ha06c,
// 16'h9c29, 16'h99f2, 16'h99cb, 16'h9bb2,
// 16'h9fa8, 16'ha58d, 16'had48, 16'hb6b4,
// 16'hc195, 16'hcdc2, 16'hdaec, 16'he8de,
// 16'hf73f, 16'h05d7, 16'h144a, 16'h2256,
// 16'h2fb0, 16'h3c12, 16'h473d, 16'h50f6,
// 16'h590b, 16'h5f53, 16'h63a9, 16'h6601,
// 16'h663e, 16'h6474, 16'h6096, 16'h5aca,
// 16'h5325, 16'h49ce, 16'h3eff, 16'h32e0,
// 16'h25c2, 16'h17d9, 16'h0979, 16'hfae4,
// 16'hec6e, 16'hde59, 16'hd0f7, 16'hc485,
// 16'hb949, 16'haf7f, 16'ha74e, 16'ha0f6,
// 16'h9c7f, 16'h9a12, 16'h99b9, 16'h9b67,
// 16'h9f2e, 16'ha4de, 16'hac71, 16'hb5ae,
// 16'hc071, 16'hcc7d, 16'hd990, 16'he773,
// 16'hf5cc, 16'h0462, 16'h12da, 16'h20f7,
// 16'h2e62, 16'h3ae4, 16'h462e, 16'h500f,
// 16'h5851, 16'h5ec7, 16'h6352, 16'h65dc,
// 16'h6651, 16'h64b8, 16'h6111, 16'h5b74,
// 16'h53fc, 16'h4ad2, 16'h4020, 16'h3426,
// 16'h271a, 16'h1944, 16'h0aee, 16'hfc58,
// 16'heddd, 16'hdfbb, 16'hd244, 16'hc5b6,
// 16'hba5a, 16'hb065, 16'ha80f, 16'ha180,
// 16'h9cdc, 16'h9a38, 16'h99a8, 16'h9b27,
// 16'h9eb5, 16'ha437, 16'hab9b, 16'hb4af,
// 16'hbf4e, 16'hcb3a, 16'hd83a, 16'he606,
// 16'hf45b, 16'h02ec, 16'h116a, 16'h1f94,
// 16'h2d16, 16'h39ae, 16'h451f, 16'h4f24,
// 16'h578f, 16'h5e3a, 16'h62f3, 16'h65b4,
// 16'h665d, 16'h64f7, 16'h6188, 16'h5c17,
// 16'h54d2, 16'h4bcd, 16'h4142, 16'h3567,
// 16'h2871, 16'h1aad, 16'h0c61, 16'hfdce,
// 16'hef4d, 16'he120, 16'hd38f, 16'hc6ef,
// 16'hbb6a, 16'hb155, 16'ha8d0, 16'ha211,
// 16'h9d3d, 16'h9a65, 16'h999c, 16'h9aec,
// 16'h9e3f, 16'ha398, 16'haac7, 16'hb3b5,
// 16'hbe2e, 16'hc9fb, 16'hd6e4, 16'he49c,
// 16'hf2e9, 16'h0176, 16'h0ffa, 16'h1e31,
// 16'h2bc3, 16'h387c, 16'h4404, 16'h4e39,
// 16'h56ca, 16'h5da5, 16'h6292, 16'h6582,
// 16'h6666, 16'h6533, 16'h61f6, 16'h5cb9,
// 16'h55a0, 16'h4cc6, 16'h4262, 16'h36a2,
// 16'h29c8, 16'h1c17, 16'h0dd0, 16'hff46,
// 16'hf0bd, 16'he282, 16'hd4e8, 16'hc81d,
// 16'hbc8b, 16'hb23d, 16'ha99d, 16'ha2a4,
// 16'h9da5, 16'h9a92, 16'h999d, 16'h9aaf,
// 16'h9dd5, 16'ha2f9, 16'ha9f8, 16'hb2c1,
// 16'hbd0f, 16'hc8c1, 16'hd58d, 16'he337,
// 16'hf176, 16'h2020, 16'h0e8a, 16'h1cc8,
// 16'h2a75, 16'h373e, 16'h42f0, 16'h4d41,
// 16'h5606, 16'h5d08, 16'h622d, 16'h654c,
// 16'h6669, 16'h6569, 16'h625e, 16'h5d59,
// 16'h5668, 16'h4dbc, 16'h437e, 16'h37d9,
// 16'h2b1f, 16'h1d7c, 16'h0f41, 16'h20be,
// 16'hf22c, 16'he3ec, 16'hd637, 16'hc95d,
// 16'hbd9f, 16'hb33a, 16'haa60, 16'ha346,
// 16'h9e0c, 16'h9aca, 16'h999e, 16'h9a7a,
// 16'h9d6f, 16'ha25e, 16'ha931, 16'hb1cc,
// 16'hbbf8, 16'hc786, 16'hd43d, 16'he1ce,
// 16'hf007, 16'hfe89, 16'h0d19, 16'h1b62,
// 16'h291d, 16'h3605, 16'h41d2, 16'h4c4b,
// 16'h5538, 16'h5c6b, 16'h61bd, 16'h6517,
// 16'h6663, 16'h659a, 16'h62c6, 16'h5dec,
// 16'h5730, 16'h4eae, 16'h4492, 16'h3916,
// 16'h2c6d, 16'h1ee1, 16'h10b4, 16'h0230,
// 16'hf3a1, 16'he553, 16'hd78e, 16'hca9a,
// 16'hbebd, 16'hb433, 16'hab2e, 16'ha3ea,
// 16'h9e77, 16'h9b0a, 16'h99a2, 16'h9a4d,
// 16'h9d0c, 16'ha1c8, 16'ha86e, 16'hb0de,
// 16'hbae0, 16'hc654, 16'hd2e8, 16'he06d,
// 16'hee95, 16'hfd13, 16'h0ba8, 16'h19f8,
// 16'h27c7, 16'h34c6, 16'h40b0, 16'h4b53,
// 16'h5465, 16'h5bc8, 16'h614c, 16'h64d7,
// 16'h665a, 16'h65c7, 16'h6324, 16'h5e80,
// 16'h57f2, 16'h4f99, 16'h45a8, 16'h3a48,
// 16'h2dbe, 16'h2043, 16'h1226, 16'h03a3,
// 16'hf517, 16'he6b9, 16'hd8e8, 16'hcbd8,
// 16'hbfe1, 16'hb52e, 16'hac04, 16'ha48d,
// 16'h9eec, 16'h9b4c, 16'h99ab, 16'h9a27,
// 16'h9cad, 16'ha138, 16'ha7b0, 16'haff2,
// 16'hb9cf, 16'hc520, 16'hd199, 16'hdf0d,
// 16'hed23, 16'hfba1, 16'h0a31, 16'h1890,
// 16'h266e, 16'h3383, 16'h3f90, 16'h4a50,
// 16'h5392, 16'h5b1f, 16'h60d6, 16'h6494,
// 16'h664a, 16'h65ee, 16'h637f, 16'h5f0e,
// 16'h58ae, 16'h5082, 16'h46b8, 16'h3b79,
// 16'h2f0c, 16'h21a5, 16'h1392, 16'h051d,
// 16'hf685, 16'he829, 16'hda3d, 16'hcd20,
// 16'hc101, 16'hb632, 16'hacdc, 16'ha534,
// 16'h9f6b, 16'h9b8c, 16'h99c0, 16'h9a03,
// 16'h9c52, 16'ha0b1, 16'ha6f2, 16'haf0b,
// 16'hb8c4, 16'hc3ec, 16'hd052, 16'hdda8,
// 16'hebb7, 16'hfa2b, 16'h08bd, 16'h1726,
// 16'h2511, 16'h3241, 16'h3e68, 16'h494f,
// 16'h52b6, 16'h5a73, 16'h6059, 16'h644d,
// 16'h6636, 16'h660e, 16'h63d5, 16'h5f96,
// 16'h5967, 16'h5168, 16'h47c3, 16'h3ca8,
// 16'h3055, 16'h2307, 16'h14ff, 16'h0693,
// 16'hf7f8, 16'he996, 16'hdb98, 16'hce67,
// 16'hc228, 16'hb738, 16'hadb5, 16'ha5e8,
// 16'h9fe5, 16'h9bdb, 16'h99d4, 16'h99e6,
// 16'h9bfe, 16'ha02c, 16'ha63b, 16'hae2a,
// 16'hb7b7, 16'hc2c3, 16'hcf03, 16'hdc4f,
// 16'hea46, 16'hf8b6, 16'h074c, 16'h15b5,
// 16'h23b7, 16'h30f9, 16'h3d3f, 16'h4847,
// 16'h51d9, 16'h59c1, 16'h5fd8, 16'h63ff,
// 16'h661c, 16'h662b, 16'h6425, 16'h6019,
// 16'h5a1c, 16'h5247, 16'h48cd, 16'h3dd2,
// 16'h319e, 16'h2463, 16'h1670, 16'h0803,
// 16'hf971, 16'heafe, 16'hdcfa, 16'hcfac,
// 16'hc356, 16'hb83e, 16'hae98, 16'ha69a,
// 16'ha068, 16'h9c2e, 16'h99ee, 16'h99cd,
// 16'h9bb2, 16'h9fa8, 16'ha58c, 16'had4a,
// 16'hb6b2, 16'hc196, 16'hcdc3, 16'hdaea,
// 16'he8df, 16'hf73f, 16'h05d8, 16'h1447,
// 16'h225a, 16'h2fac, 16'h3c15, 16'h473b,
// 16'h50f7, 16'h590b, 16'h5f52, 16'h63ac,
// 16'h65fd, 16'h6642, 16'h6471, 16'h6097,
// 16'h5acb, 16'h5323, 16'h49d2, 16'h3efa,
// 16'h32e4, 16'h25bf, 16'h17da, 16'h097a,
// 16'hfae3, 16'hec6f, 16'hde58, 16'hd0f7,
// 16'hc485, 16'hb94a, 16'haf7d, 16'ha751,
// 16'ha0f3, 16'h9c81, 16'h9a12, 16'h99b6,
// 16'h9b6b, 16'h9f2b, 16'ha4e0, 16'hac70,
// 16'hb5af, 16'hc070, 16'hcc7d, 16'hd991,
// 16'he772, 16'hf5ce, 16'h0460, 16'h12dc,
// 16'h20f4, 16'h2e66, 16'h3ae1, 16'h462f,
// 16'h500f, 16'h5852, 16'h5ec4, 16'h6357,
// 16'h65d6, 16'h6655, 16'h64b7, 16'h6110,
// 16'h5b76, 16'h53fa, 16'h4ad2, 16'h4022,
// 16'h3424, 16'h271b, 16'h1944, 16'h0aec,
// 16'hfc5b, 16'heddb, 16'hdfbd, 16'hd241,
// 16'hc5b9, 16'hba58, 16'hb066, 16'ha810,
// 16'ha17e, 16'h9cde, 16'h9a37, 16'h99a8,
// 16'h9b28, 16'h9eb3, 16'ha43a, 16'hab98,
// 16'hb4b2, 16'hbf4b, 16'hcb3c, 16'hd839,
// 16'he606, 16'hf45c, 16'h02ea, 16'h116b,
// 16'h1f95, 16'h2d14, 16'h39b1, 16'h451c,
// 16'h4f24, 16'h5792, 16'h5e36, 16'h62f8,
// 16'h65ae, 16'h6661, 16'h64f7, 16'h6186,
// 16'h5c1a, 16'h54ce, 16'h4bcf, 16'h4143,
// 16'h3565, 16'h2873, 16'h1aad, 16'h0c5f,
// 16'hfdd0, 16'hef4c, 16'he11f, 16'hd392,
// 16'hc6eb, 16'hbb6f, 16'hb151, 16'ha8d2,
// 16'ha210, 16'h9d3e, 16'h9a62, 16'h99a2,
// 16'h9ae5, 16'h9e47, 16'ha390, 16'haacc,
// 16'hb3b3, 16'hbe2e, 16'hc9fd, 16'hd6e1,
// 16'he49f, 16'hf2e7, 16'h0176, 16'h0ffa,
// 16'h1e31, 16'h2bc5, 16'h3878, 16'h4409,
// 16'h4e33, 16'h56cf, 16'h5da3, 16'h6291,
// 16'h6586, 16'h6660, 16'h6539, 16'h61f1,
// 16'h5cbd, 16'h559d, 16'h4cc9, 16'h425f,
// 16'h36a4, 16'h29c8, 16'h1c15, 16'h0dd2,
// 16'hff45, 16'hf0bd, 16'he284, 16'hd4e5,
// 16'hc821, 16'hbc86, 16'hb243, 16'ha996,
// 16'ha2ab, 16'h9da0, 16'h9a96, 16'h999a,
// 16'h9ab0, 16'h9dd5, 16'ha2f9, 16'ha9f8,
// 16'hb2c0, 16'hbd10, 16'hc8c0, 16'hd58f,
// 16'he335, 16'hf177, 16'hffff, 16'h0e8a,
// 16'h1cca, 16'h2a72, 16'h3742, 16'h42ec,
// 16'h4d44, 16'h5604, 16'h5d09, 16'h622c,
// 16'h654e, 16'h6668, 16'h6568, 16'h6261,
// 16'h5d55, 16'h566b, 16'h4dbc, 16'h437b,
// 16'h37dd, 16'h2b1c, 16'h1d7d, 16'h0f43,
// 16'h20ba, 16'hf22f, 16'he3ea, 16'hd638,
// 16'hc95e, 16'hbd9e, 16'hb339, 16'haa62,
// 16'ha345, 16'h9e0b, 16'h9acd, 16'h9999,
// 16'h9a7f, 16'h9d6c, 16'ha25f, 16'ha931,
// 16'hb1cc, 16'hbbf8, 16'hc786, 16'hd43c,
// 16'he1d0, 16'hf005, 16'hfe8b, 16'h0d17,
// 16'h1b63, 16'h291d, 16'h3604, 16'h41d4,
// 16'h4c48, 16'h553b, 16'h5c68, 16'h61c0,
// 16'h6516, 16'h6661, 16'h659d, 16'h62c2,
// 16'h5df0, 16'h572e, 16'h4eae, 16'h4493,
// 16'h3913, 16'h2c71, 16'h1edd, 16'h10b8,
// 16'h022d, 16'hf3a3, 16'he551, 16'hd78e,
// 16'hca9c, 16'hbebc, 16'hb433, 16'hab2f,
// 16'ha3e7, 16'h9e7a, 16'h9b09, 16'h99a1,
// 16'h9a4f, 16'h9d0a, 16'ha1c9, 16'ha86f,
// 16'hb0dc, 16'hbae3, 16'hc650, 16'hd2ec,
// 16'he06b, 16'hee95, 16'hfd15, 16'h0ba4,
// 16'h19fc, 16'h27c5, 16'h34c6, 16'h40b2,
// 16'h4b50, 16'h5466, 16'h5bc9, 16'h614a,
// 16'h64db, 16'h6656, 16'h65ca, 16'h6321,
// 16'h5e83, 16'h57ef, 16'h4f9c, 16'h45a6,
// 16'h3a48, 16'h2dbf, 16'h2043, 16'h1225,
// 16'h03a5, 16'hf514, 16'he6bc, 16'hd8e5,
// 16'hcbdc, 16'hbfdd, 16'hb531, 16'hac03,
// 16'ha48c, 16'h9eee, 16'h9b4a, 16'h99ad,
// 16'h9a26, 16'h9cad, 16'ha139, 16'ha7af,
// 16'haff2, 16'hb9cf, 16'hc520, 16'hd19b,
// 16'hdf0b, 16'hed24, 16'hfba0, 16'h0a32,
// 16'h1890, 16'h266c, 16'h3386, 16'h3f8d,
// 16'h4a54, 16'h538d, 16'h5b23, 16'h60d3,
// 16'h6495, 16'h664c, 16'h65ea, 16'h6383,
// 16'h5f0b, 16'h58b0, 16'h5081, 16'h46b8,
// 16'h3b7a, 16'h2f0b, 16'h21a6, 16'h1391,
// 16'h051d, 16'hf687, 16'he826, 16'hda40,
// 16'hcd1e, 16'hc102, 16'hb633, 16'hacd8,
// 16'ha539, 16'h9f67, 16'h9b8e, 16'h99c2,
// 16'h99fe, 16'h9c58, 16'ha0ab, 16'ha6f6,
// 16'haf0b, 16'hb8c1, 16'hc3f1, 16'hd04d,
// 16'hddab, 16'hebb6, 16'hfa2a, 16'h08c0,
// 16'h1723, 16'h2513, 16'h323e, 16'h3e6b,
// 16'h494c, 16'h52b9, 16'h5a72, 16'h6058,
// 16'h644e, 16'h6634, 16'h6610, 16'h63d5,
// 16'h5f96, 16'h5966, 16'h5169, 16'h47c2,
// 16'h3ca8, 16'h3057, 16'h2303, 16'h1504,
// 16'h068e, 16'hf7fc, 16'he992, 16'hdb9c,
// 16'hce63, 16'hc22c, 16'hb735, 16'hadb6,
// 16'ha5e9, 16'h9fe2, 16'h9bdf, 16'h99d2,
// 16'h99e5, 16'h9c02, 16'ha025, 16'ha642,
// 16'hae26, 16'hb7b9, 16'hc2c1, 16'hcf06,
// 16'hdc4b, 16'hea4a, 16'hf8b4, 16'h074b,
// 16'h15b7, 16'h23b6, 16'h30f9, 16'h3d40,
// 16'h4845, 16'h51db, 16'h59bf, 16'h5fdb,
// 16'h63fc, 16'h661e, 16'h662b, 16'h6423,
// 16'h601d, 16'h5a17, 16'h524b, 16'h48ca,
// 16'h3dd5, 16'h319c, 16'h2464, 16'h166e,
// 16'h0804, 16'hf973, 16'heafb, 16'hdcfe,
// 16'hcfa7, 16'hc35b, 16'hb83b, 16'hae99,
// 16'ha699, 16'ha06a, 16'h9c2c, 16'h99f1,
// 16'h99c9, 16'h9bb5, 16'h9fa6, 16'ha58e,
// 16'had49, 16'hb6b1, 16'hc199, 16'hcdbe,
// 16'hdaf1, 16'he8d8, 16'hf744, 16'h05d4,
// 16'h144b, 16'h2256, 16'h2fb0, 16'h3c12,
// 16'h473c, 16'h50f8, 16'h5909, 16'h5f54,
// 16'h63a9, 16'h6601, 16'h663e, 16'h6474,
// 16'h6096, 16'h5ac9, 16'h5326, 16'h49d0,
// 16'h3efa, 16'h32e6, 16'h25bc, 16'h17dd,
// 16'h0977, 16'hfae5, 16'hec6d, 16'hde5b,
// 16'hd0f4, 16'hc487, 16'hb948, 16'haf7f,
// 16'ha74f, 16'ha0f6, 16'h9c7c, 16'h9a17,
// 16'h99b3, 16'h9b6d, 16'h9f2a, 16'ha4e1,
// 16'hac6e, 16'hb5b0, 16'hc071, 16'hcc7b,
// 16'hd995, 16'he76e, 16'hf5cf, 16'h0460,
// 16'h12dc, 16'h20f5, 16'h2e65, 16'h3ae1,
// 16'h4630, 16'h500e, 16'h5851, 16'h5ec7,
// 16'h6353, 16'h65da, 16'h6653, 16'h64b7,
// 16'h6110, 16'h5b76, 16'h53fa, 16'h4ad3,
// 16'h4020, 16'h3426, 16'h271a, 16'h1944,
// 16'h0aec, 16'hfc5b, 16'heddc, 16'hdfbb,
// 16'hd243, 16'hc5b7, 16'hba5a, 16'hb066,
// 16'ha80e, 16'ha180, 16'h9cdc, 16'h9a39,
// 16'h99a7, 16'h9b28, 16'h9eb3, 16'ha43a,
// 16'hab97, 16'hb4b3, 16'hbf4a, 16'hcb3e,
// 16'hd837, 16'he608, 16'hf459, 16'h02ec,
// 16'h116c, 16'h1f93, 16'h2d15, 16'h39b1,
// 16'h451a, 16'h4f28, 16'h578e, 16'h5e39,
// 16'h62f5, 16'h65b1, 16'h665f, 16'h64f7,
// 16'h6186, 16'h5c1b, 16'h54ce, 16'h4bd0,
// 16'h4140, 16'h3567, 16'h2873, 16'h1aac,
// 16'h0c61, 16'hfdce, 16'hef4d, 16'he11f,
// 16'hd391, 16'hc6ec, 16'hbb6e, 16'hb152,
// 16'ha8d0, 16'ha213, 16'h9d3b, 16'h9a65,
// 16'h999f, 16'h9ae6, 16'h9e46, 16'ha393,
// 16'haac9, 16'hb3b5, 16'hbe2d, 16'hc9fc,
// 16'hd6e3, 16'he49d, 16'hf2e9, 16'h0174,
// 16'h0ffd, 16'h1e2e, 16'h2bc6, 16'h3878,
// 16'h4408, 16'h4e36, 16'h56cc, 16'h5da5,
// 16'h628f, 16'h6586, 16'h6663, 16'h6535,
// 16'h61f5, 16'h5cba, 16'h559f, 16'h4cc6,
// 16'h4263, 16'h36a0, 16'h29cc, 16'h1c11,
// 16'h0dd6, 16'hff42, 16'hf0bf, 16'he283,
// 16'hd4e2, 16'hc827, 16'hbc81, 16'hb246,
// 16'ha996, 16'ha2a8, 16'h9da3, 16'h9a94,
// 16'h999b, 16'h9ab0, 16'h9dd6, 16'ha2f6,
// 16'ha9fb, 16'hb2bf, 16'hbd0f, 16'hc8c3,
// 16'hd58a, 16'he33a, 16'hf173, 16'h2002,
// 16'h0e89, 16'h1cca, 16'h2a73, 16'h373e,
// 16'h42f1, 16'h4d41, 16'h5606, 16'h5d09,
// 16'h622a, 16'h6550, 16'h6666, 16'h656b,
// 16'h625e, 16'h5d59, 16'h5666, 16'h4dc0,
// 16'h4378, 16'h37e0, 16'h2b1a, 16'h1d7e,
// 16'h0f42, 16'h20bb, 16'hf22e, 16'he3ec,
// 16'hd635, 16'hc961, 16'hbd9c, 16'hb33a,
// 16'haa61, 16'ha345, 16'h9e0b, 16'h9ace,
// 16'h9998, 16'h9a7f, 16'h9d6d, 16'ha25d,
// 16'ha934, 16'hb1c9, 16'hbbf9, 16'hc788,
// 16'hd439, 16'he1d4, 16'hf001, 16'hfe8d,
// 16'h0d17, 16'h1b61, 16'h2921, 16'h3620,
// 16'h41d6, 16'h4c49, 16'h5538, 16'h5c6b,
// 16'h61be, 16'h6517, 16'h6662, 16'h659b,
// 16'h62c4, 16'h5def, 16'h572e, 16'h4eaf,
// 16'h4492, 16'h3915, 16'h2c6e, 16'h1ee0,
// 16'h10b5, 16'h0230, 16'hf3a2, 16'he551,
// 16'hd78f, 16'hca99, 16'hbebe, 16'hb433,
// 16'hab2e, 16'ha3ea, 16'h9e76, 16'h9b0b,
// 16'h999f, 16'h9a51, 16'h9d0a, 16'ha1c8,
// 16'ha86f, 16'hb0db, 16'hbae4, 16'hc651,
// 16'hd2ea, 16'he06d, 16'hee94, 16'hfd14,
// 16'h0ba8, 16'h19f7, 16'h27c8, 16'h34c5,
// 16'h40b2, 16'h4b51, 16'h5465, 16'h5bc9,
// 16'h614b, 16'h64d9, 16'h6659, 16'h65c5,
// 16'h6327, 16'h5e7e, 16'h57f3, 16'h4f99,
// 16'h45a8, 16'h3a47, 16'h2dbe, 16'h2045,
// 16'h1223, 16'h03a7, 16'hf513, 16'he6bc,
// 16'hd8e5, 16'hcbdc, 16'hbfde, 16'hb52f,
// 16'hac04, 16'ha48c, 16'h9eee, 16'h9b4b,
// 16'h99ab, 16'h9a27, 16'h9cad, 16'ha138,
// 16'ha7b1, 16'haff0, 16'hb9d1, 16'hc51e,
// 16'hd19c, 16'hdf09, 16'hed28, 16'hfb9c,
// 16'h0a35, 16'h188d, 16'h266e, 16'h3386,
// 16'h3f8d, 16'h4a52, 16'h5391, 16'h5b1e,
// 16'h60d8, 16'h6491, 16'h664e, 16'h65ea,
// 16'h6382, 16'h5f0c, 16'h58ae, 16'h5084,
// 16'h46b6, 16'h3b7a, 16'h2f0b, 16'h21a6,
// 16'h1392, 16'h051c, 16'hf687, 16'he826,
// 16'hda41, 16'hcd1c, 16'hc106, 16'hb62d,
// 16'hacde, 16'ha536, 16'h9f67, 16'h9b90,
// 16'h99bf, 16'h9a01, 16'h9c56, 16'ha0ac,
// 16'ha6f7, 16'haf08, 16'hb8c5, 16'hc3ec,
// 16'hd051, 16'hddaa, 16'hebb5, 16'hfa2c,
// 16'h08bc, 16'h1728, 16'h250e, 16'h3244,
// 16'h3e65, 16'h4951, 16'h52b4, 16'h5a76,
// 16'h6057, 16'h644e, 16'h6634, 16'h660f,
// 16'h63d6, 16'h5f94, 16'h596b, 16'h5163,
// 16'h47c6, 16'h3ca7, 16'h3056, 16'h2305,
// 16'h1503, 16'h068d, 16'hf7ff, 16'he98f,
// 16'hdb9e, 16'hce62, 16'hc22d, 16'hb733,
// 16'hadb9, 16'ha5e5, 16'h9fe7, 16'h9bda,
// 16'h99d6, 16'h99e3, 16'h9c20, 16'ha02b,
// 16'ha63c, 16'hae29, 16'hb7b8, 16'hc2c1,
// 16'hcf07, 16'hdc4b, 16'hea48, 16'hf8b6,
// 16'h074a, 16'h15b8, 16'h23b5, 16'h30f9,
// 16'h3d40, 16'h4846, 16'h51da, 16'h59c0,
// 16'h5fd9, 16'h63fe, 16'h661d, 16'h662b,
// 16'h6425, 16'h6019, 16'h5a1d, 16'h5244,
// 16'h48d1, 16'h3dcf, 16'h31a0, 16'h2463,
// 16'h166e, 16'h0805, 16'hf970, 16'heafe,
// 16'hdcfb, 16'hcfaa, 16'hc358, 16'hb83e,
// 16'hae97, 16'ha699, 16'ha06b, 16'h9c29,
// 16'h99f4, 16'h99c8, 16'h9bb5, 16'h9fa6,
// 16'ha58e, 16'had49, 16'hb6b2, 16'hc197,
// 16'hcdc0, 16'hdaee, 16'he8dd, 16'hf740,
// 16'h05d6, 16'h144a, 16'h2257, 16'h2faf,
// 16'h3c13, 16'h473c, 16'h50f6, 16'h590d,
// 16'h5f50, 16'h63ad, 16'h65fd, 16'h6641,
// 16'h6472, 16'h6097, 16'h5aca, 16'h5325,
// 16'h49cf, 16'h3efe, 16'h32e1, 16'h25c0,
// 16'h17db, 16'h0977, 16'hfae7, 16'hec6b,
// 16'hde5c, 16'hd0f4, 16'hc486, 16'hb94a,
// 16'haf7c, 16'ha753, 16'ha0f1, 16'h9c82,
// 16'h9a11, 16'h99b8, 16'h9b69, 16'h9f2c,
// 16'ha4e0, 16'hac70, 16'hb5ae, 16'hc072,
// 16'hcc7a, 16'hd995, 16'he76f, 16'hf5cf,
// 16'h0460, 16'h12da, 16'h20f8, 16'h2e62,
// 16'h3ae4, 16'h462e, 16'h500f, 16'h5851,
// 16'h5ec7, 16'h6352, 16'h65dc, 16'h6651,
// 16'h64b9, 16'h610f, 16'h5b76, 16'h53fb,
// 16'h4ad2, 16'h4020, 16'h3427, 16'h2717,
// 16'h1949, 16'h0ae8, 16'hfc5d, 16'hedda,
// 16'hdfbe, 16'hd23f, 16'hc5bb, 16'hba56,
// 16'hb068, 16'ha80e, 16'ha180, 16'h9cdb,
// 16'h9a3a, 16'h99a6, 16'h9b29, 16'h9eb3,
// 16'ha439, 16'hab9a, 16'hb4af, 16'hbf4e,
// 16'hcb3b, 16'hd839, 16'he607, 16'hf45a,
// 16'h02eb, 16'h116c, 16'h1f94, 16'h2d14,
// 16'h39b0, 16'h451d, 16'h4f24, 16'h5792,
// 16'h5e36, 16'h62f6, 16'h65b0, 16'h6661,
// 16'h64f5, 16'h6189, 16'h5c16, 16'h54d2,
// 16'h4bcd, 16'h4144, 16'h3564, 16'h2873,
// 16'h1aac, 16'h0c61, 16'hfdcf, 16'hef4c,
// 16'he120, 16'hd38f, 16'hc6ef, 16'hbb6b,
// 16'hb154, 16'ha8cf, 16'ha214, 16'h9d3a,
// 16'h9a66, 16'h999e, 16'h9ae8, 16'h9e44,
// 16'ha394, 16'haac9, 16'hb3b5, 16'hbe2d,
// 16'hc9fc, 16'hd6e3, 16'he49d, 16'hf2ea,
// 16'h0172, 16'h0ffe, 16'h1e2e, 16'h2bc5,
// 16'h387b, 16'h4405, 16'h4e37, 16'h56cc,
// 16'h5da4, 16'h6292, 16'h6583, 16'h6665,
// 16'h6533, 16'h61f7, 16'h5cb8, 16'h55a1,
// 16'h4cc6, 16'h4260, 16'h36a5, 16'h29c6,
// 16'h1c17, 16'h0dd1, 16'hff45, 16'hf0bd,
// 16'he285, 16'hd4e2, 16'hc824, 16'hbc84,
// 16'hb244, 16'ha997, 16'ha2a8, 16'h9da2,
// 16'h9a95, 16'h999b, 16'h9ab0, 16'h9dd4,
// 16'ha2f8, 16'ha9fb, 16'hb2be, 16'hbd11,
// 16'hc8c0, 16'hd58c, 16'he339, 16'hf174,
// 16'h2002, 16'h0e88, 16'h1ccb, 16'h2a71,
// 16'h3741, 16'h42ee, 16'h4d43, 16'h5604,
// 16'h5d0b, 16'h6228, 16'h6551, 16'h6666,
// 16'h656a, 16'h6260, 16'h5d55, 16'h566b,
// 16'h4dbb, 16'h437c, 16'h37dd, 16'h2b1c,
// 16'h1d7c, 16'h0f45, 16'h20b7, 16'hf233,
// 16'he3e6, 16'hd63b, 16'hc95b, 16'hbda1,
// 16'hb338, 16'haa61, 16'ha347, 16'h9e08,
// 16'h9acf, 16'h9999, 16'h9a7f, 16'h9d6d,
// 16'ha25c, 16'ha935, 16'hb1c7, 16'hbbfd,
// 16'hc784, 16'hd43c, 16'he1d1, 16'hf003,
// 16'hfe8c, 16'h0d18, 16'h1b61, 16'h2920,
// 16'h3601, 16'h41d5, 16'h4c49, 16'h5539,
// 16'h5c6b, 16'h61bd, 16'h6517, 16'h6662,
// 16'h659b, 16'h62c6, 16'h5deb, 16'h5731,
// 16'h4ead, 16'h4493, 16'h3915, 16'h2c6d,
// 16'h1ee1, 16'h10b4, 16'h0231, 16'hf3a1,
// 16'he552, 16'hd78c, 16'hca9e, 16'hbeba,
// 16'hb435, 16'hab2f, 16'ha3e5, 16'h9e7d,
// 16'h9b04, 16'h99a6, 16'h9a4c, 16'h9d0c,
// 16'ha1c7, 16'ha870, 16'hb0db, 16'hbae4,
// 16'hc651, 16'hd2e8, 16'he070, 16'hee91,
// 16'hfd18, 16'h0ba3, 16'h19fc, 16'h27c4,
// 16'h34c8, 16'h40b0, 16'h4b52, 16'h5465,
// 16'h5bc9, 16'h614c, 16'h64d7, 16'h665a,
// 16'h65c7, 16'h6323, 16'h5e82, 16'h57ef,
// 16'h4f9c, 16'h45a6, 16'h3a49, 16'h2dbc,
// 16'h2045, 16'h1225, 16'h03a3, 16'hf518,
// 16'he6b7, 16'hd8e9, 16'hcbd9, 16'hbfe0,
// 16'hb52e, 16'hac05, 16'ha48b, 16'h9eef,
// 16'h9b49, 16'h99ad, 16'h9a26, 16'h9cad,
// 16'ha139, 16'ha7af, 16'haff1, 16'hb9d1,
// 16'hc51e, 16'hd19c, 16'hdf0a, 16'hed25,
// 16'hfb9f, 16'h0a34, 16'h188d, 16'h2670,
// 16'h3381, 16'h3f92, 16'h4a50, 16'h5390,
// 16'h5b21, 16'h60d4, 16'h6495, 16'h664a,
// 16'h65ee, 16'h637e, 16'h5f0f, 16'h58ad,
// 16'h5084, 16'h46b6, 16'h3b7a, 16'h2f0b,
// 16'h21a5, 16'h1395, 16'h0519, 16'hf689,
// 16'he825, 16'hda40, 16'hcd1f, 16'hc102,
// 16'hb632, 16'hacda, 16'ha536, 16'h9f6a,
// 16'h9b8c, 16'h99c3, 16'h99fe, 16'h9c57,
// 16'ha0ac, 16'ha6f7, 16'haf08, 16'hb8c5,
// 16'hc3ec, 16'hd051, 16'hddaa, 16'hebb5,
// 16'hfa2c, 16'h08bd, 16'h1725, 16'h2513,
// 16'h323e, 16'h3e6a, 16'h494e, 16'h52b7,
// 16'h5a73, 16'h6058, 16'h644d, 16'h6636,
// 16'h660f, 16'h63d5, 16'h5f96, 16'h5965,
// 16'h516b, 16'h47bf, 16'h3cac, 16'h3054,
// 16'h2304, 16'h1504, 16'h068d, 16'hf7fe,
// 16'he990, 16'hdb9d, 16'hce63, 16'hc22b,
// 16'hb737, 16'hadb5, 16'ha5e7, 16'h9fe6,
// 16'h9bda, 16'h99d7, 16'h99e2, 16'h9c02,
// 16'ha028, 16'ha63e, 16'hae28, 16'hb7b9,
// 16'hc2c0, 16'hcf08, 16'hdc4a, 16'hea48,
// 16'hf8b7, 16'h0749, 16'h15b8, 16'h23b6,
// 16'h30f7, 16'h3d42, 16'h4844, 16'h51dc,
// 16'h59be, 16'h5fdc, 16'h63fa, 16'h6621,
// 16'h6627, 16'h6428, 16'h6018, 16'h5a1c,
// 16'h5247, 16'h48cd, 16'h3dd2, 16'h319e,
// 16'h2464, 16'h166d, 16'h0806, 16'hf96f,
// 16'heaff, 16'hdcfb, 16'hcfa9, 16'hc35a,
// 16'hb83a, 16'hae9c, 16'ha696, 16'ha06d,
// 16'h9c28, 16'h99f4, 16'h99c7, 16'h9bb7,
// 16'h9fa5, 16'ha58e, 16'had48, 16'hb6b3,
// 16'hc197, 16'hcdc0, 16'hdaee, 16'he8dc,
// 16'hf740, 16'h05d9, 16'h1446, 16'h2259,
// 16'h2faf, 16'h3c11, 16'h4740, 16'h50f3,
// 16'h590d, 16'h5f52, 16'h63a9, 16'h6602,
// 16'h663e, 16'h6473, 16'h6097, 16'h5aca,
// 16'h5324, 16'h49d0, 16'h3efc, 16'h32e3,
// 16'h25bf, 16'h17dc, 16'h0975, 16'hfae8,
// 16'hec6b, 16'hde5b, 16'hd0f7, 16'hc482,
// 16'hb94e, 16'haf79, 16'ha755, 16'ha0f0,
// 16'h9c83, 16'h9a10, 16'h99b9, 16'h9b68,
// 16'h9f2d, 16'ha4e0, 16'hac6f, 16'hb5af,
// 16'hc071, 16'hcc7b, 16'hd994, 16'he770,
// 16'hf5ce, 16'h0460, 16'h12dc, 16'h20f4,
// 16'h2e67, 16'h3adf, 16'h4632, 16'h500c,
// 16'h5854, 16'h5ec4, 16'h6356, 16'h65d7,
// 16'h6655, 16'h64b5, 16'h6115, 16'h5b70,
// 16'h5420, 16'h4acd, 16'h4024, 16'h3425,
// 16'h2719, 16'h1946, 16'h0aeb, 16'hfc5b,
// 16'heddc, 16'hdfbb, 16'hd243, 16'hc5b7,
// 16'hba5a, 16'hb065, 16'ha80f, 16'ha181,
// 16'h9cd9, 16'h9a3d, 16'h99a3, 16'h9b2b,
// 16'h9eb1, 16'ha43b, 16'hab99, 16'hb4ae,
// 16'hbf51, 16'hcb36, 16'hd83e, 16'he603,
// 16'hf45d, 16'h02e9, 16'h116d, 16'h1f94,
// 16'h2d14, 16'h39b1, 16'h451c, 16'h4f23,
// 16'h5794, 16'h5e35, 16'h62f7, 16'h65b1,
// 16'h665d, 16'h64fa, 16'h6183, 16'h5c1c,
// 16'h54cf, 16'h4bcd, 16'h4145, 16'h3562,
// 16'h2876, 16'h1aab, 16'h0c61, 16'hfdce,
// 16'hef4e, 16'he11c, 16'hd396, 16'hc6e8,
// 16'hbb70, 16'hb151, 16'ha8d1, 16'ha211,
// 16'h9d3e, 16'h9a62, 16'h99a0, 16'h9ae8,
// 16'h9e43, 16'ha395, 16'haac8, 16'hb3b4,
// 16'hbe30, 16'hc9f9, 16'hd6e5, 16'he49c,
// 16'hf2e9, 16'h0175, 16'h0ffb, 16'h1e30,
// 16'h2bc5, 16'h3879, 16'h4408, 16'h4e34,
// 16'h56cf, 16'h5da2, 16'h6292, 16'h6585,
// 16'h6662, 16'h6537, 16'h61f2, 16'h5cbd,
// 16'h559e, 16'h4cc6, 16'h4263, 16'h36a0,
// 16'h29ca, 16'h1c16, 16'h0dd1, 16'hff45,
// 16'hf0be, 16'he282, 16'hd4e5, 16'hc823,
// 16'hbc83, 16'hb247, 16'ha993, 16'ha2ad,
// 16'h9d9d, 16'h9a98, 16'h9999, 16'h9ab1,
// 16'h9dd5, 16'ha2f7, 16'ha9fb, 16'hb2be,
// 16'hbd12, 16'hc8be, 16'hd590, 16'he334,
// 16'hf178, 16'hffff, 16'h0e8a, 16'h1ccb,
// 16'h2a70, 16'h3742, 16'h42ee, 16'h4d41,
// 16'h5607, 16'h5d07, 16'h622d, 16'h654e,
// 16'h6667, 16'h656a, 16'h625e, 16'h5d59,
// 16'h5667, 16'h4dbe, 16'h437b, 16'h37dd,
// 16'h2b1c, 16'h1d7c, 16'h0f44, 16'h20b9,
// 16'hf231, 16'he3e8, 16'hd639, 16'hc95d,
// 16'hbd9f, 16'hb339, 16'haa61, 16'ha346,
// 16'h9e0b, 16'h9acb, 16'h999d, 16'h9a7a,
// 16'h9d71, 16'ha25a, 16'ha936, 16'hb1c7,
// 16'hbbfc, 16'hc783, 16'hd43e, 16'he1cf,
// 16'hf005, 16'hfe8b, 16'h0d17, 16'h1b63,
// 16'h291d, 16'h3604, 16'h41d3, 16'h4c4a,
// 16'h553a, 16'h5c67, 16'h61c3, 16'h6511,
// 16'h6667, 16'h6598, 16'h62c6, 16'h5dec,
// 16'h5732, 16'h4eab, 16'h4495, 16'h3913,
// 16'h2c6d, 16'h1ee4, 16'h10b1, 16'h0233,
// 16'hf39e, 16'he555, 16'hd78b, 16'hca9e,
// 16'hbebb, 16'hb432, 16'hab32, 16'ha3e4,
// 16'h9e7c, 16'h9b08, 16'h99a0, 16'h9a51,
// 16'h9d08, 16'ha1cb, 16'ha86e, 16'hb0db,
// 16'hbae5, 16'hc64e, 16'hd2ed, 16'he06c,
// 16'hee93, 16'hfd16, 16'h0ba5, 16'h19fa,
// 16'h27c7, 16'h34c4, 16'h40b3, 16'h4b4f,
// 16'h5469, 16'h5bc5, 16'h614f, 16'h64d4,
// 16'h665e, 16'h65c1, 16'h632b, 16'h5e7a,
// 16'h57f6, 16'h4f97, 16'h45a8, 16'h3a49,
// 16'h2dbc, 16'h2046, 16'h1222, 16'h03a7,
// 16'hf515, 16'he6b9, 16'hd8e9, 16'hcbd7,
// 16'hbfe2, 16'hb52e, 16'hac04, 16'ha48c,
// 16'h9eee, 16'h9b49, 16'h99af, 16'h9a23,
// 16'h9cb1, 16'ha134, 16'ha7b4, 16'hafed,
// 16'hb9d3, 16'hc51f, 16'hd199, 16'hdf0e,
// 16'hed20, 16'hfba4, 16'h0a2f, 16'h1892,
// 16'h266c, 16'h3384, 16'h3f90, 16'h4a4f,
// 16'h5394, 16'h5b1d, 16'h60d7, 16'h6494,
// 16'h6649, 16'h65f0, 16'h637d, 16'h5f0f,
// 16'h58ae, 16'h5082, 16'h46b9, 16'h3b78,
// 16'h2f0b, 16'h21a7, 16'h1391, 16'h051e,
// 16'hf684, 16'he829, 16'hda3f, 16'hcd1d,
// 16'hc105, 16'hb62e, 16'hacde, 16'ha535,
// 16'h9f68, 16'h9b90, 16'h99bd, 16'h9a04,
// 16'h9c53, 16'ha0af, 16'ha6f5, 16'haf08,
// 16'hb8c6, 16'hc3ea, 16'hd055, 16'hdda5,
// 16'hebb9, 16'hfa29, 16'h08c0, 16'h1723,
// 16'h2513, 16'h323f, 16'h3e69, 16'h494f,
// 16'h52b6, 16'h5a73, 16'h6059, 16'h644c,
// 16'h6637, 16'h660e, 16'h63d5, 16'h5f96,
// 16'h5967, 16'h5168, 16'h47c2, 16'h3caa,
// 16'h3053, 16'h2308, 16'h1520, 16'h0690,
// 16'hf7fb, 16'he992, 16'hdb9c, 16'hce65,
// 16'hc229, 16'hb736, 16'hadb7, 16'ha5e6,
// 16'h9fe7, 16'h9bdb, 16'h99d3, 16'h99e6,
// 16'h9c20, 16'ha028, 16'ha640, 16'hae26,
// 16'hb7ba, 16'hc2c0, 16'hcf07, 16'hdc4b,
// 16'hea48, 16'hf8b7, 16'h0749, 16'h15b8,
// 16'h23b5, 16'h30fa, 16'h3d3d, 16'h484b,
// 16'h51d4, 16'h59c5, 16'h5fd7, 16'h63fd,
// 16'h661f, 16'h6629, 16'h6426, 16'h601a,
// 16'h5a1a, 16'h5248, 16'h48cc, 16'h3dd4,
// 16'h319c, 16'h2466, 16'h166b, 16'h0807,
// 16'hf96f, 16'heaff, 16'hdcfb, 16'hcfaa,
// 16'hc357, 16'hb83e, 16'hae98, 16'ha699,
// 16'ha06b, 16'h9c29, 16'h99f3, 16'h99c9,
// 16'h9bb4, 16'h9fa7, 16'ha58d, 16'had49,
// 16'hb6b3, 16'hc196, 16'hcdc0, 16'hdaef,
// 16'he8da, 16'hf744, 16'h05d3, 16'h144b,
// 16'h2257, 16'h2fae, 16'h3c14, 16'h473c,
// 16'h50f5, 16'h590d, 16'h5f51, 16'h63ab,
// 16'h6620, 16'h663f, 16'h6472, 16'h6098,
// 16'h5ac9, 16'h5326, 16'h49ce, 16'h3efe,
// 16'h32e1, 16'h25c2, 16'h17d8, 16'h097a,
// 16'hfae4, 16'hec6d, 16'hde5b, 16'hd0f5,
// 16'hc485, 16'hb94b, 16'haf7b, 16'ha753,
// 16'ha0f3, 16'h9c7f, 16'h9a15, 16'h99b3,
// 16'h9b6d, 16'h9f2a, 16'ha4e1, 16'hac70,
// 16'hb5ad, 16'hc073, 16'hcc79, 16'hd996,
// 16'he76d, 16'hf5d1, 16'h045e, 16'h12dc,
// 16'h20f7, 16'h2e62, 16'h3ae4, 16'h462e,
// 16'h500f, 16'h5851, 16'h5ec7, 16'h6352,
// 16'h65dd, 16'h6650, 16'h64b8, 16'h6111,
// 16'h5b74, 16'h53fd, 16'h4ad0, 16'h4022,
// 16'h3424, 16'h271c, 16'h1943, 16'h0aed,
// 16'hfc5a, 16'heddb, 16'hdfbe, 16'hd240,
// 16'hc5b9, 16'hba59, 16'hb065, 16'ha80f,
// 16'ha181, 16'h9cda, 16'h9a3b, 16'h99a5,
// 16'h9b28, 16'h9eb5, 16'ha438, 16'hab99,
// 16'hb4b1, 16'hbf4c, 16'hcb3c, 16'hd839,
// 16'he606, 16'hf45b, 16'h02eb, 16'h116c,
// 16'h1f94, 16'h2d14, 16'h39b0, 16'h451d,
// 16'h4f25, 16'h5791, 16'h5e37, 16'h62f5,
// 16'h65b2, 16'h665e, 16'h64f9, 16'h6184,
// 16'h5c1c, 16'h54cd, 16'h4bd1, 16'h4140,
// 16'h3567, 16'h2872, 16'h1aad, 16'h0c60,
// 16'hfdcf, 16'hef4c, 16'he120, 16'hd391,
// 16'hc6eb, 16'hbb6f, 16'hb150, 16'ha8d4,
// 16'ha20f, 16'h9d3d, 16'h9a65, 16'h999d,
// 16'h9aeb, 16'h9e41, 16'ha395, 16'haaca,
// 16'hb3b2, 16'hbe31, 16'hc9fa, 16'hd6e3,
// 16'he49d, 16'hf2e9, 16'h0174, 16'h0ffe,
// 16'h1e2d, 16'h2bc6, 16'h3879, 16'h4407,
// 16'h4e36, 16'h56cd, 16'h5da3, 16'h6292,
// 16'h6583, 16'h6666, 16'h6532, 16'h61f7,
// 16'h5cb8, 16'h55a2, 16'h4cc5, 16'h4261,
// 16'h36a4, 16'h29c6, 16'h1c18, 16'h0dd0,
// 16'hff45, 16'hf0bf, 16'he281, 16'hd4e6,
// 16'hc821, 16'hbc86, 16'hb243, 16'ha997,
// 16'ha2a9, 16'h9da0, 16'h9a98, 16'h9998,
// 16'h9ab2, 16'h9dd5, 16'ha2f5, 16'ha9fd,
// 16'hb2be, 16'hbd10, 16'hc8c2, 16'hd58c,
// 16'he337, 16'hf176, 16'h2020, 16'h0e89,
// 16'h1ccc, 16'h2a70, 16'h3741, 16'h42ee,
// 16'h4d44, 16'h5602, 16'h5d0d, 16'h6225,
// 16'h6555, 16'h6662, 16'h656e, 16'h625c,
// 16'h5d58, 16'h5669, 16'h4dbc, 16'h437d,
// 16'h37db, 16'h2b1e, 16'h1d7c, 16'h0f41,
// 16'h20bd, 16'hf22d, 16'he3eb, 16'hd639,
// 16'hc95a, 16'hbda3, 16'hb336, 16'haa63,
// 16'ha343, 16'h9e0e, 16'h9aca, 16'h999c,
// 16'h9a7e, 16'h9d6b, 16'ha25f, 16'ha933,
// 16'hb1c8, 16'hbbfd, 16'hc782, 16'hd43f,
// 16'he1ce, 16'hf006, 16'hfe8a, 16'h0d19,
// 16'h1b60, 16'h2921, 16'h3620, 16'h41d6,
// 16'h4c49, 16'h5538, 16'h5c6c, 16'h61bc,
// 16'h6518, 16'h6662, 16'h659a, 16'h62c6,
// 16'h5dec, 16'h5731, 16'h4ead, 16'h4493,
// 16'h3913, 16'h2c70, 16'h1edf, 16'h10b6,
// 16'h022e, 16'hf3a3, 16'he551, 16'hd78e,
// 16'hca9b, 16'hbebc, 16'hb434, 16'hab2f,
// 16'ha3e6, 16'h9e7b, 16'h9b08, 16'h99a1,
// 16'h9a50, 16'h9d09, 16'ha1c9, 16'ha870,
// 16'hb0da, 16'hbae4, 16'hc651, 16'hd2ea,
// 16'he06c, 16'hee97, 16'hfd11, 16'h0ba9,
// 16'h19f7, 16'h27c8, 16'h34c5, 16'h40b3,
// 16'h4b4f, 16'h5467, 16'h5bc8, 16'h614c,
// 16'h64d8, 16'h6658, 16'h65c8, 16'h6324,
// 16'h5e81, 16'h57f0, 16'h4f9a, 16'h45a8,
// 16'h3a47, 16'h2dbf, 16'h2043, 16'h1225,
// 16'h03a5, 16'hf514, 16'he6bc, 16'hd8e5,
// 16'hcbdc, 16'hbfde, 16'hb530, 16'hac02,
// 16'ha48e, 16'h9eed, 16'h9b4a, 16'h99ae,
// 16'h9a24, 16'h9caf, 16'ha137, 16'ha7b2,
// 16'hafed, 16'hb9d5, 16'hc51b, 16'hd19d,
// 16'hdf0c, 16'hed21, 16'hfba3, 16'h0a2f,
// 16'h1892, 16'h266c, 16'h3385, 16'h3f8f,
// 16'h4a50, 16'h5392, 16'h5b1e, 16'h60d7,
// 16'h6493, 16'h664c, 16'h65ec, 16'h6380,
// 16'h5f0d, 16'h58af, 16'h5083, 16'h46b5,
// 16'h3b7d, 16'h2f07, 16'h21a9, 16'h1392,
// 16'h0519, 16'hf68b, 16'he822, 16'hda44,
// 16'hcd1a, 16'hc106, 16'hb62f, 16'hacdc,
// 16'ha537, 16'h9f66, 16'h9b92, 16'h99bc,
// 16'h9a04, 16'h9c54, 16'ha0ad, 16'ha6f6,
// 16'haf0a, 16'hb8c2, 16'hc3ef, 16'hd04f,
// 16'hddaa, 16'hebb7, 16'hfa2a, 16'h08be,
// 16'h1724, 16'h2514, 16'h323d, 16'h3e6c,
// 16'h494c, 16'h52b6, 16'h5a76, 16'h6056,
// 16'h644e, 16'h6636, 16'h660d, 16'h63d6,
// 16'h5f96, 16'h5966, 16'h516a, 16'h47c0,
// 16'h3caa, 16'h3055, 16'h2304, 16'h1505,
// 16'h068b, 16'hf801, 16'he98c, 16'hdba1,
// 16'hce60, 16'hc22d, 16'hb735, 16'hadb7,
// 16'ha5e6, 16'h9fe6, 16'h9bda, 16'h99d7,
// 16'h99e1, 16'h9c04, 16'ha026, 16'ha640,
// 16'hae26, 16'hb7bb, 16'hc2be, 16'hcf09,
// 16'hdc49, 16'hea4a, 16'hf8b4, 16'h074e,
// 16'h15b2, 16'h23ba, 16'h30f5, 16'h3d43,
// 16'h4844, 16'h51dc, 16'h59bd, 16'h5fdc,
// 16'h63fc, 16'h661e, 16'h662a, 16'h6426,
// 16'h6019, 16'h5a1b, 16'h5248, 16'h48cb,
// 16'h3dd4, 16'h319e, 16'h2463, 16'h166f,
// 16'h0804, 16'hf970, 16'heaff, 16'hdcfa,
// 16'hcfab, 16'hc358, 16'hb83d, 16'hae98,
// 16'ha69a, 16'ha069, 16'h9c2a, 16'h99f4,
// 16'h99c7, 16'h9bb6, 16'h9fa7, 16'ha58b,
// 16'had4b, 16'hb6b2, 16'hc195, 16'hcdc3,
// 16'hdaec, 16'he8dd, 16'hf741, 16'h05d5,
// 16'h144a, 16'h2258, 16'h2fae, 16'h3c14,
// 16'h473a, 16'h50f9, 16'h5908, 16'h5f56,
// 16'h63a9, 16'h65ff, 16'h6640, 16'h6471,
// 16'h6099, 16'h5ac9, 16'h5325, 16'h49cf,
// 16'h3efd, 16'h32e2, 16'h25c1, 16'h17d8,
// 16'h097a, 16'hfae5, 16'hec6c, 16'hde5b,
// 16'hd0f5, 16'hc486, 16'hb949, 16'haf7e,
// 16'ha750, 16'ha0f4, 16'h9c7f, 16'h9a14,
// 16'h99b5, 16'h9b6c, 16'h9f2a, 16'ha4e1,
// 16'hac6f, 16'hb5af, 16'hc071, 16'hcc7b,
// 16'hd994, 16'he770, 16'hf5cd, 16'h0462,
// 16'h12d9, 16'h20f8, 16'h2e63, 16'h3ae2,
// 16'h462f, 16'h500f, 16'h5851, 16'h5ec7,
// 16'h6353, 16'h65da, 16'h6652, 16'h64b9,
// 16'h610e, 16'h5b79, 16'h53f7, 16'h4ad4,
// 16'h4021, 16'h3424, 16'h271c, 16'h1943,
// 16'h0aec, 16'hfc5c, 16'hedda, 16'hdfbd,
// 16'hd241, 16'hc5b9, 16'hba58, 16'hb068,
// 16'ha80c, 16'ha182, 16'h9cda, 16'h9a3a,
// 16'h99a8, 16'h9b27, 16'h9eb4, 16'ha438,
// 16'hab9a, 16'hb4b0, 16'hbf4e, 16'hcb3a,
// 16'hd839, 16'he607, 16'hf45b, 16'h02ea,
// 16'h116d, 16'h1f91, 16'h2d18, 16'h39af,
// 16'h451c, 16'h4f26, 16'h578e, 16'h5e3b,
// 16'h62f3, 16'h65b3, 16'h665e, 16'h64f7,
// 16'h6188, 16'h5c16, 16'h54d4, 16'h4bcb,
// 16'h4144, 16'h3566, 16'h2870, 16'h1ab0,
// 16'h0c5e, 16'hfdd0, 16'hef4c, 16'he11e,
// 16'hd394, 16'hc6ea, 16'hbb6e, 16'hb152,
// 16'ha8d1, 16'ha212, 16'h9d3c, 16'h9a64,
// 16'h999f, 16'h9ae8, 16'h9e44, 16'ha393,
// 16'haaca, 16'hb3b4, 16'hbe2e, 16'hc9fc,
// 16'hd6e1, 16'he4a0, 16'hf2e6, 16'h0177,
// 16'h0ffb, 16'h1e2f, 16'h2bc5, 16'h387a,
// 16'h4406, 16'h4e37, 16'h56cc, 16'h5da4,
// 16'h6292, 16'h6583, 16'h6664, 16'h6535,
// 16'h61f4, 16'h5cbc, 16'h559d, 16'h4cc9,
// 16'h425f, 16'h36a4, 16'h29c7, 16'h1c17,
// 16'h0dd0, 16'hff48, 16'hf0b9, 16'he288,
// 16'hd4e0, 16'hc825, 16'hbc85, 16'hb242,
// 16'ha999, 16'ha2a7, 16'h9da2, 16'h9a96,
// 16'h9999, 16'h9ab3, 16'h9dd1, 16'ha2fb,
// 16'ha9f8, 16'hb2c0, 16'hbd11, 16'hc8bf,
// 16'hd58e, 16'he337, 16'hf175, 16'h2001,
// 16'h0e8a, 16'h1cc9, 16'h2a73, 16'h3740,
// 16'h42ee, 16'h4d43, 16'h5604, 16'h5d0a,
// 16'h622a, 16'h6550, 16'h6666, 16'h6569,
// 16'h6261, 16'h5d55, 16'h566b, 16'h4dbb,
// 16'h437c, 16'h37dd, 16'h2b1d, 16'h1d7b,
// 16'h0f44, 16'h20ba, 16'hf22f, 16'he3eb,
// 16'hd636, 16'hc95f, 16'hbd9e, 16'hb339,
// 16'haa62, 16'ha344, 16'h9e0d, 16'h9aca,
// 16'h999e, 16'h9a7a, 16'h9d6f, 16'ha25d,
// 16'ha932, 16'hb1cd, 16'hbbf5, 16'hc78a,
// 16'hd439, 16'he1d1, 16'hf006, 16'hfe88,
// 16'h0d1b, 16'h1b60, 16'h291e, 16'h3606,
// 16'h41cf, 16'h4c4f, 16'h5534, 16'h5c6d,
// 16'h61bd, 16'h6518, 16'h6660, 16'h659e,
// 16'h62c0, 16'h5df3, 16'h572c, 16'h4eaf,
// 16'h4492, 16'h3914, 16'h2c70, 16'h1ede,
// 16'h10b8, 16'h022c, 16'hf3a4, 16'he551,
// 16'hd78e, 16'hca9a, 16'hbec0, 16'hb42e,
// 16'hab34, 16'ha3e4, 16'h9e7b, 16'h9b08,
// 16'h99a2, 16'h9a4e, 16'h9d0b, 16'ha1c9,
// 16'ha86e, 16'hb0dc, 16'hbae4, 16'hc64f,
// 16'hd2ec, 16'he06b, 16'hee95, 16'hfd16,
// 16'h0ba3, 16'h19fd, 16'h27c2, 16'h34c9,
// 16'h40b1, 16'h4b4f, 16'h546a, 16'h5bc3,
// 16'h6150, 16'h64d5, 16'h665b, 16'h65c7,
// 16'h6323, 16'h5e81, 16'h57f1, 16'h4f9a,
// 16'h45a7, 16'h3a48, 16'h2dbe, 16'h2045,
// 16'h1223, 16'h03a6, 16'hf513, 16'he6be,
// 16'hd8e3, 16'hcbde, 16'hbfdb, 16'hb532,
// 16'hac03, 16'ha48c, 16'h9eef, 16'h9b48,
// 16'h99ae, 16'h9a26, 16'h9cad, 16'ha138,
// 16'ha7b1, 16'hafef, 16'hb9d2, 16'hc51e,
// 16'hd19b, 16'hdf0b, 16'hed24, 16'hfba0,
// 16'h0a32, 16'h1890, 16'h266c, 16'h3386,
// 16'h3f8d, 16'h4a53, 16'h538f, 16'h5b21,
// 16'h60d5, 16'h6494, 16'h664a, 16'h65ef,
// 16'h637d, 16'h5f10, 16'h58ad, 16'h5083,
// 16'h46b8, 16'h3b78, 16'h2f0d, 16'h21a4,
// 16'h1395, 16'h0519, 16'hf689, 16'he825,
// 16'hda41, 16'hcd1d, 16'hc104, 16'hb630,
// 16'hacdb, 16'ha537, 16'h9f67, 16'h9b91,
// 16'h99bd, 16'h9a04, 16'h9c52, 16'ha0b0,
// 16'ha6f3, 16'haf0b, 16'hb8c4, 16'hc3ec,
// 16'hd051, 16'hddaa, 16'hebb4, 16'hfa2e,
// 16'h08bb, 16'h1727, 16'h2510, 16'h3241,
// 16'h3e69, 16'h494d, 16'h52b9, 16'h5a70,
// 16'h605b, 16'h644c, 16'h6635, 16'h6610,
// 16'h63d5, 16'h5f94, 16'h596a, 16'h5164,
// 16'h47c6, 16'h3ca7, 16'h3056, 16'h2305,
// 16'h1502, 16'h068f, 16'hf7fc, 16'he993,
// 16'hdb9a, 16'hce65, 16'hc22c, 16'hb732,
// 16'hadbc, 16'ha5e2, 16'h9fe8, 16'h9bdb,
// 16'h99d4, 16'h99e4, 16'h9c02, 16'ha027,
// 16'ha63f, 16'hae28, 16'hb7b7, 16'hc2c4,
// 16'hcf03, 16'hdc4e, 16'hea46, 16'hf8b8,
// 16'h0749, 16'h15b7, 16'h23b7, 16'h30f6,
// 16'h3d44, 16'h4843, 16'h51db, 16'h59bf,
// 16'h5fdb, 16'h63fc, 16'h661f, 16'h6629,
// 16'h6425, 16'h601c, 16'h5a18, 16'h5249,
// 16'h48cd, 16'h3dd0, 16'h31a2, 16'h245f,
// 16'h1673, 16'h07ff, 16'hf975, 16'heafb,
// 16'hdcfd, 16'hcfa9, 16'hc358, 16'hb83d,
// 16'hae99, 16'ha698, 16'ha06b, 16'h9c2a,
// 16'h99f2, 16'h99c9, 16'h9bb5, 16'h9fa6,
// 16'ha58e, 16'had48, 16'hb6b3, 16'hc196,
// 16'hcdc1, 16'hdaee, 16'he8da, 16'hf745,
// 16'h05d1, 16'h144e, 16'h2253, 16'h2fb3,
// 16'h3c0f, 16'h4740, 16'h50f4, 16'h590c,
// 16'h5f52, 16'h63aa, 16'h6620, 16'h6641,
// 16'h6470, 16'h6099, 16'h5ac8, 16'h5326,
// 16'h49cf, 16'h3efd, 16'h32e2, 16'h25c1,
// 16'h17d8, 16'h097a, 16'hfae5, 16'hec6c,
// 16'hde5c, 16'hd0f2, 16'hc48a, 16'hb947,
// 16'haf7e, 16'ha751, 16'ha0f2, 16'h9c82,
// 16'h9a13, 16'h99b4, 16'h9b6d, 16'h9f29,
// 16'ha4e3, 16'hac6d, 16'hb5b0, 16'hc071,
// 16'hcc7b, 16'hd995, 16'he76d, 16'hf5d1,
// 16'h045e, 16'h12dd, 16'h20f5, 16'h2e64,
// 16'h3ae3, 16'h462e, 16'h500f, 16'h5850,
// 16'h5ec9, 16'h6351, 16'h65dd, 16'h664f,
// 16'h64ba, 16'h6110, 16'h5b74, 16'h53fd,
// 16'h4acf, 16'h4024, 16'h3423, 16'h271b,
// 16'h1944, 16'h0aeb, 16'hfc5d, 16'hedda,
// 16'hdfbc, 16'hd243, 16'hc5b5, 16'hba5d,
// 16'hb063, 16'ha811, 16'ha17e, 16'h9cdc,
// 16'h9a39, 16'h99a8, 16'h9b27, 16'h9eb5,
// 16'ha437, 16'hab9b, 16'hb4ae, 16'hbf50,
// 16'hcb39, 16'hd83a, 16'he607, 16'hf459,
// 16'h02ec, 16'h116d, 16'h1f91, 16'h2d18,
// 16'h39ad, 16'h451f, 16'h4f22, 16'h5795,
// 16'h5e33, 16'h62f9, 16'h65af, 16'h665f,
// 16'h64f9, 16'h6184, 16'h5c1c, 16'h54cd,
// 16'h4bd1, 16'h413f, 16'h3569, 16'h2870,
// 16'h1aaf, 16'h0c5f, 16'hfdce, 16'hef4e,
// 16'he11e, 16'hd393, 16'hc6ea, 16'hbb6f,
// 16'hb151, 16'ha8d1, 16'ha213, 16'h9d3b,
// 16'h9a64, 16'h99a0, 16'h9ae7, 16'h9e44,
// 16'ha394, 16'haac9, 16'hb3b4, 16'hbe2f,
// 16'hc9fb, 16'hd6e2, 16'he49f, 16'hf2e7,
// 16'h0176, 16'h0ffb, 16'h1e30, 16'h2bc4,
// 16'h387a, 16'h4407, 16'h4e35, 16'h56cf,
// 16'h5da0, 16'h6296, 16'h657f, 16'h6669,
// 16'h6530, 16'h61f8, 16'h5cb9, 16'h55a0,
// 16'h4cc5, 16'h4263, 16'h36a1, 16'h29ca,
// 16'h1c15, 16'h0dd0, 16'hff47, 16'hf0bb,
// 16'he286, 16'hd4e2, 16'hc824, 16'hbc84,
// 16'hb244, 16'ha996, 16'ha2aa, 16'h9da0,
// 16'h9a97, 16'h9999, 16'h9ab2, 16'h9dd2,
// 16'ha2fb, 16'ha9f7, 16'hb2c2, 16'hbd0e,
// 16'hc8c1, 16'hd58e, 16'he336, 16'hf176,
// 16'h2020, 16'h0e8a, 16'h1cca, 16'h2a72,
// 16'h3740, 16'h42ee, 16'h4d44, 16'h5603,
// 16'h5d0a, 16'h622b, 16'h654f, 16'h6667,
// 16'h6569, 16'h625f, 16'h5d58, 16'h5668,
// 16'h4dbe, 16'h437a, 16'h37de, 16'h2b1b,
// 16'h1d7e, 16'h0f41, 16'h20bd, 16'hf22d,
// 16'he3eb, 16'hd638, 16'hc95c, 16'hbda1,
// 16'hb337, 16'haa63, 16'ha344, 16'h9e0c,
// 16'h9acb, 16'h999d, 16'h9a7b, 16'h9d6f,
// 16'ha25c, 16'ha933, 16'hb1cc, 16'hbbf7,
// 16'hc788, 16'hd43a, 16'he1d1, 16'hf005,
// 16'hfe8a, 16'h0d18, 16'h1b63, 16'h291c,
// 16'h3606, 16'h41d1, 16'h4c4b, 16'h5538,
// 16'h5c6b, 16'h61be, 16'h6517, 16'h6661,
// 16'h659c, 16'h62c3, 16'h5df0, 16'h572e,
// 16'h4eae, 16'h4493, 16'h3912, 16'h2c71,
// 16'h1edf, 16'h10b5, 16'h0230, 16'hf3a0,
// 16'he553, 16'hd78f, 16'hca98, 16'hbec0,
// 16'hb42f, 16'hab32, 16'ha3e6, 16'h9e7b,
// 16'h9b06, 16'h99a4, 16'h9a4d, 16'h9d0b,
// 16'ha1ca, 16'ha86c, 16'hb0df, 16'hbae1,
// 16'hc652, 16'hd2ea, 16'he06c, 16'hee95,
// 16'hfd15, 16'h0ba4, 16'h19fc, 16'h27c4,
// 16'h34c7, 16'h40b2, 16'h4b4f, 16'h5468,
// 16'h5bc7, 16'h614c, 16'h64d8, 16'h665a,
// 16'h65c5, 16'h6326, 16'h5e80, 16'h57f0,
// 16'h4f9c, 16'h45a5, 16'h3a49, 16'h2dbf,
// 16'h2042, 16'h1227, 16'h03a2, 16'hf517,
// 16'he6ba, 16'hd8e7, 16'hcbda, 16'hbfdf,
// 16'hb52e, 16'hac05, 16'ha48b, 16'h9ef0,
// 16'h9b47, 16'h99b0, 16'h9a23, 16'h9caf,
// 16'ha137, 16'ha7b1, 16'haff1, 16'hb9d0,
// 16'hc51f, 16'hd19b, 16'hdf0b, 16'hed25,
// 16'hfb9f, 16'h0a32, 16'h1891, 16'h266b,
// 16'h3387, 16'h3f8c, 16'h4a54, 16'h538f,
// 16'h5b20, 16'h60d6, 16'h6494, 16'h6649,
// 16'h65f1, 16'h637b, 16'h5f12, 16'h58ab,
// 16'h5084, 16'h46b7, 16'h3b79, 16'h2f0d,
// 16'h21a4, 16'h1394, 16'h051a, 16'hf688,
// 16'he826, 16'hda40, 16'hcd1e, 16'hc103,
// 16'hb631, 16'hacda, 16'ha538, 16'h9f67,
// 16'h9b90, 16'h99be, 16'h9a02, 16'h9c55,
// 16'ha0ae, 16'ha6f4, 16'haf0b, 16'hb8c2,
// 16'hc3ef, 16'hd04f, 16'hddaa, 16'hebb6,
// 16'hfa2a, 16'h08bf, 16'h1725, 16'h2510,
// 16'h3242, 16'h3e68, 16'h494c, 16'h52bb,
// 16'h5a6f, 16'h605c, 16'h644b, 16'h6635,
// 16'h6610, 16'h63d5, 16'h5f96, 16'h5966,
// 16'h5169, 16'h47c1, 16'h3cab, 16'h3054,
// 16'h2304, 16'h1505, 16'h068c, 16'hf7ff,
// 16'he98f, 16'hdb9e, 16'hce62, 16'hc22d,
// 16'hb733, 16'hadba, 16'ha5e3, 16'h9fe9,
// 16'h9bd8, 16'h99d8, 16'h99e1, 16'h9c03,
// 16'ha027, 16'ha63e, 16'hae2a, 16'hb7b6,
// 16'hc2c3, 16'hcf05, 16'hdc4c, 16'hea47,
// 16'hf8b8, 16'h0748, 16'h15b9, 16'h23b5,
// 16'h30f9, 16'h3d3f, 16'h4848, 16'h51d7,
// 16'h59c2, 16'h5fda, 16'h63fb, 16'h6620,
// 16'h6628, 16'h6427, 16'h6019, 16'h5a1b,
// 16'h5247, 16'h48cd, 16'h3dd3, 16'h319e,
// 16'h2463, 16'h166e, 16'h0805, 16'hf96f,
// 16'heb01, 16'hdcf8, 16'hcfad, 16'hc355,
// 16'hb83f, 16'hae97, 16'ha69a, 16'ha06a,
// 16'h9c2b, 16'h99f0, 16'h99cb, 16'h9bb4,
// 16'h9fa7, 16'ha58d, 16'had49, 16'hb6b1,
// 16'hc198, 16'hcdc1, 16'hdaed, 16'he8dc,
// 16'hf741, 16'h05d6, 16'h144a, 16'h2257,
// 16'h2fae, 16'h3c14, 16'h473c, 16'h50f6,
// 16'h590c, 16'h5f51, 16'h63ad, 16'h65fc,
// 16'h6643, 16'h6470, 16'h6098, 16'h5acb,
// 16'h5322, 16'h49d2, 16'h3efb, 16'h32e3,
// 16'h25c1, 16'h17d8, 16'h097b, 16'hfae1,
// 16'hec71, 16'hde58, 16'hd0f6, 16'hc487,
// 16'hb947, 16'haf7f, 16'ha751, 16'ha0f1,
// 16'h9c84, 16'h9a10, 16'h99b6, 16'h9b6c,
// 16'h9f29, 16'ha4e4, 16'hac6c, 16'hb5b1,
// 16'hc06e, 16'hcc7f, 16'hd990, 16'he774,
// 16'hf5ca, 16'h0464, 16'h12d8, 16'h20f8,
// 16'h2e63, 16'h3ae2, 16'h4630, 16'h500e,
// 16'h5851, 16'h5ec7, 16'h6353, 16'h65da,
// 16'h6654, 16'h64b4, 16'h6115, 16'h5b71,
// 16'h53ff, 16'h4acf, 16'h4022, 16'h3424,
// 16'h271d, 16'h1941, 16'h0af0, 16'hfc56,
// 16'heddf, 16'hdfbb, 16'hd241, 16'hc5bb,
// 16'hba55, 16'hb069, 16'ha80d, 16'ha181,
// 16'h9cdb, 16'h9a3a, 16'h99a6, 16'h9b29,
// 16'h9eb3, 16'ha439, 16'hab99, 16'hb4b0,
// 16'hbf4e, 16'hcb3b, 16'hd838, 16'he608,
// 16'hf459, 16'h02ec, 16'h116c, 16'h1f93,
// 16'h2d16, 16'h39ae, 16'h451e, 16'h4f24,
// 16'h5791, 16'h5e38, 16'h62f5, 16'h65b1,
// 16'h665f, 16'h64f7, 16'h6187, 16'h5c19,
// 16'h54d0, 16'h4bce, 16'h4142, 16'h3567,
// 16'h2870, 16'h1ab1, 16'h0c5b, 16'hfdd4,
// 16'hef48, 16'he122, 16'hd390, 16'hc6ed,
// 16'hbb6d, 16'hb151, 16'ha8d3, 16'ha210,
// 16'h9d3d, 16'h9a64, 16'h999e, 16'h9ae9,
// 16'h9e44, 16'ha393, 16'haac9, 16'hb3b6,
// 16'hbe2b, 16'hca20, 16'hd6de, 16'he4a1,
// 16'hf2e6, 16'h0177, 16'h0ffb, 16'h1e2f,
// 16'h2bc5, 16'h387a, 16'h4406, 16'h4e37,
// 16'h56cc, 16'h5da4, 16'h6292, 16'h6582,
// 16'h6667, 16'h6530, 16'h61fb, 16'h5cb4,
// 16'h55a4, 16'h4cc3, 16'h4264, 16'h36a1,
// 16'h29c9, 16'h1c15, 16'h0dd2, 16'hff44,
// 16'hf0c0, 16'he280, 16'hd4e6, 16'hc823,
// 16'hbc83, 16'hb246, 16'ha995, 16'ha2a9,
// 16'h9da2, 16'h9a95, 16'h999a, 16'h9ab1,
// 16'h9dd5, 16'ha2f7, 16'ha9fa, 16'hb2bf,
// 16'hbd10, 16'hc8c2, 16'hd58c, 16'he337,
// 16'hf176, 16'hffff, 16'h0e8c, 16'h1cc8,
// 16'h2a73, 16'h3741, 16'h42ec, 16'h4d45,
// 16'h5603, 16'h5d0b, 16'h6229, 16'h6550,
// 16'h6667, 16'h6568, 16'h6262, 16'h5d54,
// 16'h566b, 16'h4dbc, 16'h437b, 16'h37dd,
// 16'h2b1c, 16'h1d7d, 16'h0f42, 16'h20bb,
// 16'hf22f, 16'he3ea, 16'hd638, 16'hc95d,
// 16'hbd9f, 16'hb33a, 16'haa60, 16'ha347,
// 16'h9e09, 16'h9ace, 16'h999b, 16'h9a7d,
// 16'h9d6c, 16'ha25f, 16'ha931, 16'hb1cd,
// 16'hbbf7, 16'hc787, 16'hd43a, 16'he1d3,
// 16'hf002, 16'hfe8d, 16'h0d16, 16'h1b64,
// 16'h291b, 16'h3607, 16'h41d1, 16'h4c4a,
// 16'h553b, 16'h5c66, 16'h61c3, 16'h6513,
// 16'h6664, 16'h659a, 16'h62c4, 16'h5df0,
// 16'h572d, 16'h4eb0, 16'h4491, 16'h3915,
// 16'h2c6d, 16'h1ee2, 16'h10b4, 16'h0231,
// 16'hf3a0, 16'he553, 16'hd78c, 16'hca9d,
// 16'hbebc, 16'hb432, 16'hab31, 16'ha3e6,
// 16'h9e7a, 16'h9b09, 16'h999f, 16'h9a52,
// 16'h9d08, 16'ha1cb, 16'ha86d, 16'hb0dc,
// 16'hbae4, 16'hc650, 16'hd2eb, 16'he06b,
// 16'hee97, 16'hfd11, 16'h0baa, 16'h19f6,
// 16'h27c8, 16'h34c5, 16'h40b2, 16'h4b50,
// 16'h5468, 16'h5bc6, 16'h614d, 16'h64d8,
// 16'h6658, 16'h65c8, 16'h6324, 16'h5e80,
// 16'h57f2, 16'h4f9a, 16'h45a6, 16'h3a49,
// 16'h2dbd, 16'h2045, 16'h1224, 16'h03a6,
// 16'hf513, 16'he6bd, 16'hd8e3, 16'hcbde,
// 16'hbfdd, 16'hb52f, 16'hac05, 16'ha48a,
// 16'h9ef1, 16'h9b46, 16'h99b0, 16'h9a24,
// 16'h9caf, 16'ha138, 16'ha7af, 16'haff1,
// 16'hb9d1, 16'hc520, 16'hd198, 16'hdf0f,
// 16'hed20, 16'hfba3, 16'h0a31, 16'h188f,
// 16'h266e, 16'h3383, 16'h3f90, 16'h4a51,
// 16'h5390, 16'h5b21, 16'h60d3, 16'h6497,
// 16'h6648, 16'h65ef, 16'h637f, 16'h5f0c,
// 16'h58b1, 16'h5080, 16'h46b9, 16'h3b7a,
// 16'h2f09, 16'h21a8, 16'h1391, 16'h051c,
// 16'hf688, 16'he825, 16'hda40, 16'hcd1f,
// 16'hc102, 16'hb631, 16'hacda, 16'ha537,
// 16'h9f69, 16'h9b8e, 16'h99bf, 16'h9a02,
// 16'h9c54, 16'ha0b0, 16'ha6f2, 16'haf0c,
// 16'hb8c3, 16'hc3ee, 16'hd04f, 16'hddab,
// 16'hebb4, 16'hfa2d, 16'h08be, 16'h1722,
// 16'h2516, 16'h323b, 16'h3e6e, 16'h494a,
// 16'h52b9, 16'h5a72, 16'h6059, 16'h644d,
// 16'h6635, 16'h6610, 16'h63d3, 16'h5f98,
// 16'h5965, 16'h5169, 16'h47c3, 16'h3ca8,
// 16'h3056, 16'h2304, 16'h1503, 16'h068e,
// 16'hf7fe, 16'he990, 16'hdb9d, 16'hce63,
// 16'hc22b, 16'hb736, 16'hadb6, 16'ha5e7,
// 16'h9fe6, 16'h9bdb, 16'h99d4, 16'h99e5,
// 16'h9bff, 16'ha02b, 16'ha63d, 16'hae27,
// 16'hb7ba, 16'hc2bf, 16'hcf09, 16'hdc49,
// 16'hea49, 16'hf8b6, 16'h074b, 16'h15b5,
// 16'h23b8, 16'h30f7, 16'h3d41, 16'h4847,
// 16'h51d7, 16'h59c3, 16'h5fd7, 16'h63ff,
// 16'h661d, 16'h662a, 16'h6425, 16'h601b,
// 16'h5a19, 16'h524a, 16'h48c9, 16'h3dd6,
// 16'h319b, 16'h2466, 16'h166d, 16'h0804,
// 16'hf971, 16'heafe, 16'hdcfb, 16'hcfab,
// 16'hc356, 16'hb83e, 16'hae99, 16'ha698,
// 16'ha06c, 16'h9c28, 16'h99f4, 16'h99c9,
// 16'h9bb4, 16'h9fa6, 16'ha58f, 16'had47,
// 16'hb6b4, 16'hc196, 16'hcdc1, 16'hdaed,
// 16'he8dd, 16'hf740, 16'h05d6, 16'h144b,
// 16'h2256, 16'h2fb0, 16'h3c12, 16'h473c,
// 16'h50f8, 16'h590a, 16'h5f52, 16'h63ad,
// 16'h65fb, 16'h6645, 16'h646e, 16'h6099,
// 16'h5aca, 16'h5324, 16'h49d1, 16'h3efa,
// 16'h32e5, 16'h25bd, 16'h17de, 16'h0975,
// 16'hfae7, 16'hec6c, 16'hde5a, 16'hd0f6,
// 16'hc485, 16'hb94a, 16'haf7c, 16'ha753,
// 16'ha0f1, 16'h9c82, 16'h9a11, 16'h99b7,
// 16'h9b6b, 16'h9f2a, 16'ha4e1, 16'hac6f,
// 16'hb5af, 16'hc072, 16'hcc7a, 16'hd993,
// 16'he772, 16'hf5cb, 16'h0464, 16'h12d8,
// 16'h20f8, 16'h2e62, 16'h3ae4, 16'h462e,
// 16'h500f, 16'h5852, 16'h5ec4, 16'h6357,
// 16'h65d7, 16'h6655, 16'h64b6, 16'h6111,
// 16'h5b75, 16'h53fc, 16'h4ad1, 16'h4021,
// 16'h3425, 16'h271b, 16'h1943, 16'h0aee,
// 16'hfc58, 16'hedde, 16'hdfba, 16'hd245,
// 16'hc5b4, 16'hba5c, 16'hb064, 16'ha810,
// 16'ha180, 16'h9cdb, 16'h9a39, 16'h99a7,
// 16'h9b29, 16'h9eb2, 16'ha43b, 16'hab96,
// 16'hb4b4, 16'hbf4a, 16'hcb3d, 16'hd839,
// 16'he605, 16'hf45d, 16'h02e9, 16'h116c,
// 16'h1f95, 16'h2d13, 16'h39b2, 16'h451b,
// 16'h4f25, 16'h5791, 16'h5e37, 16'h62f6,
// 16'h65b1, 16'h665e, 16'h64f8, 16'h6186,
// 16'h5c1a, 16'h54cf, 16'h4bcf, 16'h4141,
// 16'h3567, 16'h2872, 16'h1aac, 16'h0c63,
// 16'hfdcb, 16'hef51, 16'he11a, 16'hd396,
// 16'hc6e8, 16'hbb71, 16'hb150, 16'ha8d2,
// 16'ha211, 16'h9d3c, 16'h9a64, 16'h99a1,
// 16'h9ae5, 16'h9e46, 16'ha393, 16'haac9,
// 16'hb3b5, 16'hbe2d, 16'hc9fd, 16'hd6e1,
// 16'he49f, 16'hf2e7, 16'h0176, 16'h0ffc,
// 16'h1e2e, 16'h2bc6, 16'h3879, 16'h4407,
// 16'h4e36, 16'h56cc, 16'h5da5, 16'h6290,
// 16'h6586, 16'h6662, 16'h6536, 16'h61f3,
// 16'h5cbd, 16'h559c, 16'h4cca, 16'h425e,
// 16'h36a5, 16'h29c7, 16'h1c16, 16'h0dd2,
// 16'hff44, 16'hf0be, 16'he283, 16'hd4e5,
// 16'hc822, 16'hbc84, 16'hb246, 16'ha993,
// 16'ha2ad, 16'h9d9f, 16'h9a95, 16'h999c,
// 16'h9aaf, 16'h9dd6, 16'ha2f7, 16'ha9fa,
// 16'hb2c0, 16'hbd0e, 16'hc8c4, 16'hd58a,
// 16'he339, 16'hf175, 16'hffff, 16'h0e8c,
// 16'h1cc8, 16'h2a73, 16'h3741, 16'h42ed,
// 16'h4d44, 16'h5603, 16'h5d0a, 16'h622b,
// 16'h654f, 16'h6667, 16'h6569, 16'h6260,
// 16'h5d55, 16'h566c, 16'h4db9, 16'h437f,
// 16'h37da, 16'h2b1e, 16'h1d7b, 16'h0f44,
// 16'h20ba, 16'hf22f, 16'he3ea, 16'hd638,
// 16'hc95d, 16'hbda0, 16'hb338, 16'haa62,
// 16'ha345, 16'h9e0b, 16'h9acd, 16'h9999,
// 16'h9a81, 16'h9d69, 16'ha261, 16'ha930,
// 16'hb1cc, 16'hbbf8, 16'hc788, 16'hd43a,
// 16'he1d1, 16'hf004, 16'hfe8b, 16'h0d18,
// 16'h1b63, 16'h291d, 16'h3604, 16'h41d1,
// 16'h4c4d, 16'h5537, 16'h5c6b, 16'h61bf,
// 16'h6514, 16'h6664, 16'h659b, 16'h62c4,
// 16'h5dee, 16'h5730, 16'h4ead, 16'h4492,
// 16'h3916, 16'h2c6d, 16'h1ee1, 16'h10b5,
// 16'h022f, 16'hf3a2, 16'he552, 16'hd78d,
// 16'hca9b, 16'hbebe, 16'hb431, 16'hab31,
// 16'ha3e6, 16'h9e79, 16'h9b0a, 16'h99a0,
// 16'h9a50, 16'h9d0a, 16'ha1c8, 16'ha870,
// 16'hb0db, 16'hbae3, 16'hc651, 16'hd2ea,
// 16'he06d, 16'hee95, 16'hfd13, 16'h0ba7,
// 16'h19f9, 16'h27c6, 16'h34c7, 16'h40b1,
// 16'h4b50, 16'h5468, 16'h5bc6, 16'h614d,
// 16'h64d7, 16'h665a, 16'h65c6, 16'h6326,
// 16'h5e7e, 16'h57f3, 16'h4f98, 16'h45aa,
// 16'h3a45, 16'h2dc0, 16'h2043, 16'h1225,
// 16'h03a5, 16'hf514, 16'he6bc, 16'hd8e4,
// 16'hcbde, 16'hbfdb, 16'hb533, 16'hac20,
// 16'ha48f, 16'h9eec, 16'h9b4b, 16'h99ad,
// 16'h9a25, 16'h9cae, 16'ha138, 16'ha7b0,
// 16'haff1, 16'hb9d0, 16'hc51f, 16'hd19b,
// 16'hdf0c, 16'hed22, 16'hfba2, 16'h0a30,
// 16'h1892, 16'h266b, 16'h3386, 16'h3f8d,
// 16'h4a53, 16'h538f, 16'h5b22, 16'h60d3,
// 16'h6496, 16'h6649, 16'h65ee, 16'h637f,
// 16'h5f0e, 16'h58ae, 16'h5083, 16'h46b7,
// 16'h3b7a, 16'h2f0a, 16'h21a7, 16'h1392,
// 16'h051c, 16'hf687, 16'he826, 16'hda41,
// 16'hcd1b, 16'hc107, 16'hb62d, 16'hacde,
// 16'ha535, 16'h9f68, 16'h9b8f, 16'h99c0,
// 16'h9a01, 16'h9c55, 16'ha0ae, 16'ha6f4,
// 16'haf0b, 16'hb8c3, 16'hc3ed, 16'hd052,
// 16'hdda7, 16'hebb8, 16'hfa2a, 16'h08be,
// 16'h1725, 16'h2511, 16'h3240, 16'h3e6a,
// 16'h494d, 16'h52b8, 16'h5a71, 16'h605b,
// 16'h644a, 16'h6639, 16'h660c, 16'h63d7,
// 16'h5f94, 16'h5969, 16'h5166, 16'h47c4,
// 16'h3ca8, 16'h3055, 16'h2306, 16'h1502,
// 16'h068f, 16'hf7fb, 16'he993, 16'hdb9b,
// 16'hce64, 16'hc22c, 16'hb733, 16'hadb9,
// 16'ha5e5, 16'h9fe7, 16'h9bda, 16'h99d5,
// 16'h99e4, 16'h9c01, 16'ha029, 16'ha63d,
// 16'hae29, 16'hb7b8, 16'hc2c0, 16'hcf09,
// 16'hdc48, 16'hea4b, 16'hf8b4, 16'h074b,
// 16'h15b7, 16'h23b6, 16'h30f9, 16'h3d3f,
// 16'h4847, 16'h51d9, 16'h59c1, 16'h5fd9,
// 16'h63fd, 16'h661e, 16'h6629, 16'h6428,
// 16'h6017, 16'h5a1c, 16'h5247, 16'h48cc,
// 16'h3dd4, 16'h319e, 16'h2461, 16'h1672,
// 16'h0820, 16'hf974, 16'heafc, 16'hdcfd,
// 16'hcfa8, 16'hc359, 16'hb83d, 16'hae97,
// 16'ha69c, 16'ha067, 16'h9c2d, 16'h99f0,
// 16'h99cb, 16'h9bb3, 16'h9fa8, 16'ha58c,
// 16'had4a, 16'hb6b1, 16'hc199, 16'hcdbd,
// 16'hdaf2, 16'he8d7, 16'hf746, 16'h05d2,
// 16'h144c, 16'h2256, 16'h2faf, 16'h3c13,
// 16'h473c, 16'h50f7, 16'h590b, 16'h5f52,
// 16'h63ab, 16'h65fe, 16'h6642, 16'h6470,
// 16'h6099, 16'h5ac9, 16'h5324, 16'h49d1,
// 16'h3efa, 16'h32e6, 16'h25bc, 16'h17de,
// 16'h0975, 16'hfae6, 16'hec6f, 16'hde56,
// 16'hd0fa, 16'hc482, 16'hb94c, 16'haf7b,
// 16'ha754, 16'ha0f0, 16'h9c82, 16'h9a13,
// 16'h99b4, 16'h9b6e, 16'h9f28, 16'ha4e2,
// 16'hac6f, 16'hb5ae, 16'hc072, 16'hcc7c,
// 16'hd991, 16'he772, 16'hf5cd, 16'h0460,
// 16'h12dd, 16'h20f4, 16'h2e65, 16'h3ae2,
// 16'h462e, 16'h5010, 16'h5850, 16'h5ec9,
// 16'h6351, 16'h65dc, 16'h6650, 16'h64ba,
// 16'h610f, 16'h5b77, 16'h53f9, 16'h4ad4,
// 16'h401f, 16'h3426, 16'h271b, 16'h1943,
// 16'h0aee, 16'hfc59, 16'heddd, 16'hdfba,
// 16'hd245, 16'hc5b5, 16'hba5b, 16'hb064,
// 16'ha810, 16'ha180, 16'h9cda, 16'h9a3b,
// 16'h99a5, 16'h9b29, 16'h9eb4, 16'ha438,
// 16'hab9a, 16'hb4af, 16'hbf4f, 16'hcb39,
// 16'hd83b, 16'he606, 16'hf45a, 16'h02ec,
// 16'h116a, 16'h1f96, 16'h2d12, 16'h39b3,
// 16'h451b, 16'h4f24, 16'h5793, 16'h5e34,
// 16'h62f8, 16'h65b0, 16'h6660, 16'h64f7,
// 16'h6186, 16'h5c1a, 16'h54ce, 16'h4bd1,
// 16'h4140, 16'h3567, 16'h2871, 16'h1ab0,
// 16'h0c5d, 16'hfdd1, 16'hef4b, 16'he11e,
// 16'hd395, 16'hc6e9, 16'hbb6e, 16'hb153,
// 16'ha8cf, 16'ha214, 16'h9d3a, 16'h9a66,
// 16'h999d, 16'h9aea, 16'h9e42, 16'ha395,
// 16'haac9, 16'hb3b3, 16'hbe30, 16'hc9fa,
// 16'hd6e4, 16'he49c, 16'hf2e9, 16'h0175,
// 16'h0ffc, 16'h1e2f, 16'h2bc5, 16'h3879,
// 16'h4407, 16'h4e37, 16'h56cc, 16'h5da3,
// 16'h6293, 16'h6582, 16'h6666, 16'h6533,
// 16'h61f5, 16'h5cbb, 16'h559e, 16'h4cc9,
// 16'h425e, 16'h36a5, 16'h29c7, 16'h1c16,
// 16'h0dd2, 16'hff44, 16'hf0be, 16'he284,
// 16'hd4e3, 16'hc824, 16'hbc83, 16'hb244,
// 16'ha998, 16'ha2a8, 16'h9da2, 16'h9a95,
// 16'h9999, 16'h9ab2, 16'h9dd4, 16'ha2f8,
// 16'ha9fa, 16'hb2c0, 16'hbd0d, 16'hc8c6,
// 16'hd587, 16'he33c, 16'hf173, 16'h2001,
// 16'h0e8b, 16'h1cc7, 16'h2a76, 16'h373c,
// 16'h42f3, 16'h4d3e, 16'h5609, 16'h5d05,
// 16'h622f, 16'h654c, 16'h6667, 16'h656c,
// 16'h625c, 16'h5d5a, 16'h5667, 16'h4dbd,
// 16'h437c, 16'h37dc, 16'h2b1d, 16'h1d7c,
// 16'h0f43, 16'h20bb, 16'hf22e, 16'he3eb,
// 16'hd637, 16'hc95d, 16'hbda0, 16'hb339,
// 16'haa60, 16'ha347, 16'h9e09, 16'h9ace,
// 16'h999b, 16'h9a7d, 16'h9d6c, 16'ha260,
// 16'ha92f, 16'hb1cf, 16'hbbf5, 16'hc789,
// 16'hd439, 16'he1d3, 16'hf002, 16'hfe8d,
// 16'h0d16, 16'h1b63, 16'h291e, 16'h3604,
// 16'h41d2, 16'h4c4b, 16'h5538, 16'h5c6a,
// 16'h61c0, 16'h6514, 16'h6664, 16'h659a,
// 16'h62c4, 16'h5def, 16'h572e, 16'h4eaf,
// 16'h4492, 16'h3914, 16'h2c6e, 16'h1ee2,
// 16'h10b2, 16'h0233, 16'hf39e, 16'he555,
// 16'hd78b, 16'hca9d, 16'hbebb, 16'hb434,
// 16'hab2f, 16'ha3e7, 16'h9e7a, 16'h9b08,
// 16'h99a1, 16'h9a50, 16'h9d09, 16'ha1cb,
// 16'ha86c, 16'hb0df, 16'hbadf, 16'hc655,
// 16'hd2e6, 16'he071, 16'hee91, 16'hfd17,
// 16'h0ba4, 16'h19fa, 16'h27c7, 16'h34c5,
// 16'h40b3, 16'h4b4f, 16'h5467, 16'h5bc8,
// 16'h614c, 16'h64d8, 16'h6659, 16'h65c6,
// 16'h6327, 16'h5e7d, 16'h57f5, 16'h4f97,
// 16'h45a8, 16'h3a49, 16'h2dbd, 16'h2045,
// 16'h1224, 16'h03a4, 16'hf516, 16'he6ba,
// 16'hd8e7, 16'hcbdb, 16'hbfdd, 16'hb530,
// 16'hac03, 16'ha48d, 16'h9eef, 16'h9b48,
// 16'h99ad, 16'h9a27, 16'h9cac, 16'ha13a,
// 16'ha7ae, 16'haff2, 16'hb9d0, 16'hc520,
// 16'hd19a, 16'hdf0b, 16'hed25, 16'hfb9f,
// 16'h0a33, 16'h188f, 16'h266d, 16'h3385,
// 16'h3f8f, 16'h4a50, 16'h5392, 16'h5b1f,
// 16'h60d6, 16'h6494, 16'h664a, 16'h65ee,
// 16'h637e, 16'h5f10, 16'h58ac, 16'h5085,
// 16'h46b5, 16'h3b7a, 16'h2f0c, 16'h21a4,
// 16'h1395, 16'h051a, 16'hf687, 16'he827,
// 16'hda3f, 16'hcd1f, 16'hc102, 16'hb632,
// 16'hacd9, 16'ha53a, 16'h9f64, 16'h9b92,
// 16'h99bd, 16'h9a03, 16'h9c54, 16'ha0af,
// 16'ha6f2, 16'haf0e, 16'hb8bf, 16'hc3f1,
// 16'hd04f, 16'hddaa, 16'hebb5, 16'hfa2c,
// 16'h08be, 16'h1724, 16'h2513, 16'h323f,
// 16'h3e68, 16'h4951, 16'h52b3, 16'h5a76,
// 16'h6058, 16'h644c, 16'h6636, 16'h660f,
// 16'h63d4, 16'h5f98, 16'h5965, 16'h5169,
// 16'h47c2, 16'h3ca9, 16'h3055, 16'h2305,
// 16'h1503, 16'h068e, 16'hf7fd, 16'he990,
// 16'hdb9f, 16'hce60, 16'hc22f, 16'hb732,
// 16'hadb9, 16'ha5e6, 16'h9fe5, 16'h9bdc,
// 16'h99d4, 16'h99e5, 16'h9c20, 16'ha029,
// 16'ha63e, 16'hae27, 16'hb7ba, 16'hc2c0,
// 16'hcf07, 16'hdc4b, 16'hea48, 16'hf8b6,
// 16'h074b, 16'h15b6, 16'h23b7, 16'h30f7,
// 16'h3d42, 16'h4845, 16'h51d9, 16'h59c3,
// 16'h5fd5, 16'h6402, 16'h6619, 16'h662f,
// 16'h6421, 16'h601e, 16'h5a16, 16'h524c,
// 16'h48c9, 16'h3dd6, 16'h319b, 16'h2466,
// 16'h166d, 16'h0805, 16'hf970, 16'heaff,
// 16'hdcfa, 16'hcfab, 16'hc357, 16'hb83f,
// 16'hae95, 16'ha69d, 16'ha066, 16'h9c2e,
// 16'h99f0, 16'h99c9, 16'h9bb6, 16'h9fa5,
// 16'ha58e, 16'had49, 16'hb6b1, 16'hc198,
// 16'hcdc1, 16'hdaec, 16'he8dd, 16'hf741,
// 16'h05d4, 16'h144e, 16'h2252, 16'h2fb3,
// 16'h3c11, 16'h473d, 16'h50f6, 16'h590b,
// 16'h5f52, 16'h63ac, 16'h65fe, 16'h6642,
// 16'h646f, 16'h609a, 16'h5ac7, 16'h5326,
// 16'h49d1, 16'h3efa, 16'h32e5, 16'h25bd,
// 16'h17dc, 16'h0978, 16'hfae5, 16'hec6d,
// 16'hde5a, 16'hd0f5, 16'hc488, 16'hb946,
// 16'haf80, 16'ha750, 16'ha0f3, 16'h9c81,
// 16'h9a12, 16'h99b6, 16'h9b6b, 16'h9f2c,
// 16'ha4de, 16'hac72, 16'hb5ac, 16'hc074,
// 16'hcc7a, 16'hd993, 16'he770, 16'hf5cf,
// 16'h045e, 16'h12df, 16'h20f2, 16'h2e67,
// 16'h3ae0, 16'h4630, 16'h500e, 16'h5852,
// 16'h5ec6, 16'h6354, 16'h65d9, 16'h6653,
// 16'h64b7, 16'h6112, 16'h5b74, 16'h53fb,
// 16'h4ad2, 16'h4020, 16'h3427, 16'h2719,
// 16'h1945, 16'h0aec, 16'hfc59, 16'hedde,
// 16'hdfba, 16'hd244, 16'hc5b7, 16'hba58,
// 16'hb067, 16'ha80f, 16'ha17e, 16'h9cdf,
// 16'h9a35, 16'h99aa, 16'h9b27, 16'h9eb3,
// 16'ha43a, 16'hab98, 16'hb4b0, 16'hbf4f,
// 16'hcb39, 16'hd83b, 16'he605, 16'hf45c,
// 16'h02e9, 16'h116e, 16'h1f91, 16'h2d18,
// 16'h39ae, 16'h451d, 16'h4f24, 16'h5791,
// 16'h5e38, 16'h62f5, 16'h65b2, 16'h665d,
// 16'h64f9, 16'h6185, 16'h5c1a, 16'h54d1,
// 16'h4bcb, 16'h4146, 16'h3562, 16'h2875,
// 16'h1aac, 16'h0c60, 16'hfdd0, 16'hef4b,
// 16'he120, 16'hd391, 16'hc6ec, 16'hbb6e,
// 16'hb152, 16'ha8d1, 16'ha211, 16'h9d3d,
// 16'h9a64, 16'h999e, 16'h9aea, 16'h9e41,
// 16'ha397, 16'haac6, 16'hb3b8, 16'hbe2a,
// 16'hc9ff, 16'hd6e0, 16'he49f, 16'hf2e9,
// 16'h0173, 16'h0fff, 16'h1e2b, 16'h2bc8,
// 16'h3878, 16'h4408, 16'h4e36, 16'h56cc,
// 16'h5da3, 16'h6293, 16'h6583, 16'h6665,
// 16'h6534, 16'h61f3, 16'h5cbe, 16'h559c,
// 16'h4cc9, 16'h4260, 16'h36a2, 16'h29ca,
// 16'h1c14, 16'h0dd4, 16'hff42, 16'hf0c0,
// 16'he281, 16'hd4e7, 16'hc81f, 16'hbc89,
// 16'hb240, 16'ha998, 16'ha2aa, 16'h9d9f,
// 16'h9a98, 16'h9999, 16'h9aaf, 16'h9dd8,
// 16'ha2f4, 16'ha9fd, 16'hb2bd, 16'hbd12,
// 16'hc8bf, 16'hd58f, 16'he335, 16'hf177,
// 16'h2020, 16'h0e88, 16'h1ccd, 16'h2a70,
// 16'h3741, 16'h42f0, 16'h4d3e, 16'h560a,
// 16'h5d05, 16'h622e, 16'h654d, 16'h6667,
// 16'h656a, 16'h6260, 16'h5d56, 16'h566a,
// 16'h4dba, 16'h437e, 16'h37dc, 16'h2b1c,
// 16'h1d7e, 16'h0f41, 16'h20bc, 16'hf22e,
// 16'he3ea, 16'hd638, 16'hc95e, 16'hbd9e,
// 16'hb33a, 16'haa60, 16'ha347, 16'h9e09,
// 16'h9acf, 16'h9998, 16'h9a80, 16'h9d6b,
// 16'ha25f, 16'ha933, 16'hb1c9, 16'hbbfb,
// 16'hc783, 16'hd440, 16'he1cb, 16'hf00a,
// 16'hfe86, 16'h0d1b, 16'h1b61, 16'h291e,
// 16'h3604, 16'h41d2, 16'h4c4b, 16'h5539,
// 16'h5c69, 16'h61c0, 16'h6515, 16'h6663,
// 16'h659a, 16'h62c6, 16'h5dec, 16'h5731,
// 16'h4ead, 16'h4493, 16'h3913, 16'h2c70,
// 16'h1edf, 16'h10b5, 16'h0232, 16'hf39d,
// 16'he557, 16'hd789, 16'hca9e, 16'hbebc,
// 16'hb432, 16'hab31, 16'ha3e5, 16'h9e7b,
// 16'h9b08, 16'h99a2, 16'h9a4e, 16'h9d0c,
// 16'ha1c7, 16'ha870, 16'hb0db, 16'hbae3,
// 16'hc652, 16'hd2e8, 16'he070, 16'hee90,
// 16'hfd19, 16'h0ba2, 16'h19fc, 16'h27c5,
// 16'h34c7, 16'h40b1, 16'h4b50, 16'h5468,
// 16'h5bc5, 16'h6150, 16'h64d5, 16'h665a,
// 16'h65c7, 16'h6324, 16'h5e80, 16'h57f2,
// 16'h4f9a, 16'h45a5, 16'h3a4c, 16'h2db9,
// 16'h2049, 16'h1220, 16'h03a9, 16'hf511,
// 16'he6be, 16'hd8e4, 16'hcbdc, 16'hbfdf,
// 16'hb52e, 16'hac05, 16'ha48b, 16'h9eef,
// 16'h9b49, 16'h99ae, 16'h9a25, 16'h9cad,
// 16'ha139, 16'ha7b0, 16'haff0, 16'hb9d2,
// 16'hc51d, 16'hd19c, 16'hdf0c, 16'hed22,
// 16'hfba2, 16'h0a30, 16'h1892, 16'h266b,
// 16'h3386, 16'h3f8e, 16'h4a51, 16'h5392,
// 16'h5b1d, 16'h60d8, 16'h6493, 16'h664c,
// 16'h65eb, 16'h6381, 16'h5f0c, 16'h58b0,
// 16'h5083, 16'h46b5, 16'h3b7c, 16'h2f09,
// 16'h21a7, 16'h1392, 16'h051c, 16'hf687,
// 16'he827, 16'hda3e, 16'hcd1f, 16'hc104,
// 16'hb62e, 16'hacde, 16'ha534, 16'h9f69,
// 16'h9b90, 16'h99be, 16'h9a01, 16'h9c57,
// 16'ha0aa, 16'ha6f8, 16'haf09, 16'hb8c3,
// 16'hc3ef, 16'hd04e, 16'hddab, 16'hebb6,
// 16'hfa2a, 16'h08c0, 16'h1721, 16'h2516,
// 16'h323c, 16'h3e6c, 16'h494c, 16'h52b8,
// 16'h5a72, 16'h605a, 16'h644a, 16'h6639,
// 16'h660d, 16'h63d5, 16'h5f97, 16'h5965,
// 16'h5169, 16'h47c4, 16'h3ca6, 16'h3058,
// 16'h2302, 16'h1505, 16'h068e, 16'hf7fc,
// 16'he992, 16'hdb9b, 16'hce65, 16'hc22b,
// 16'hb734, 16'hadb9, 16'ha5e4, 16'h9fe9,
// 16'h9bd8, 16'h99d7, 16'h99e2, 16'h9c03,
// 16'ha027, 16'ha640, 16'hae25, 16'hb7bb,
// 16'hc2bf, 16'hcf08, 16'hdc4a, 16'hea49,
// 16'hf8b6, 16'h074a, 16'h15b7, 16'h23b6,
// 16'h30f8, 16'h3d40, 16'h4848, 16'h51d8,
// 16'h59c1, 16'h5fd9, 16'h63fd, 16'h661e,
// 16'h662a, 16'h6426, 16'h6018, 16'h5a1e,
// 16'h5244, 16'h48ce, 16'h3dd3, 16'h319e,
// 16'h2462, 16'h1671, 16'h0820, 16'hf974,
// 16'heafd, 16'hdcfb, 16'hcfab, 16'hc356,
// 16'hb83f, 16'hae96, 16'ha69c, 16'ha067,
// 16'h9c2d, 16'h99f1, 16'h99ca, 16'h9bb3,
// 16'h9fa8, 16'ha58b, 16'had4c, 16'hb6b0,
// 16'hc198, 16'hcdc0, 16'hdaed, 16'he8dd,
// 16'hf741, 16'h05d5, 16'h144b, 16'h2254,
// 16'h2fb3, 16'h3c0f, 16'h4740, 16'h50f3,
// 16'h590d, 16'h5f52, 16'h63aa, 16'h6620,
// 16'h6640, 16'h6471, 16'h6099, 16'h5ac8,
// 16'h5326, 16'h49cf, 16'h3efd, 16'h32e2,
// 16'h25c1, 16'h17d8, 16'h097b, 16'hfae3,
// 16'hec6e, 16'hde5a, 16'hd0f5, 16'hc487,
// 16'hb948, 16'haf7e, 16'ha751, 16'ha0f3,
// 16'h9c81, 16'h9a11, 16'h99b7, 16'h9b6b,
// 16'h9f2b, 16'ha4e1, 16'hac6e, 16'hb5b0,
// 16'hc070, 16'hcc7d, 16'hd991, 16'he772,
// 16'hf5ce, 16'h045f, 16'h12de, 16'h20f2,
// 16'h2e67, 16'h3ae1, 16'h462f, 16'h5010,
// 16'h584f, 16'h5ec8, 16'h6353, 16'h65db,
// 16'h6651, 16'h64b9, 16'h610e, 16'h5b78,
// 16'h53f9, 16'h4ad3, 16'h4020, 16'h3426,
// 16'h2719, 16'h1946, 16'h0aea, 16'hfc5c,
// 16'heddc, 16'hdfbb, 16'hd243, 16'hc5b6,
// 16'hba5a, 16'hb067, 16'ha80d, 16'ha182,
// 16'h9cd9, 16'h9a3a, 16'h99a8, 16'h9b26,
// 16'h9eb6, 16'ha437, 16'hab9a, 16'hb4b0,
// 16'hbf4e, 16'hcb3a, 16'hd839, 16'he608,
// 16'hf459, 16'h02ed, 16'h116a, 16'h1f94,
// 16'h2d16, 16'h39ae, 16'h451f, 16'h4f22,
// 16'h5793, 16'h5e37, 16'h62f4, 16'h65b3,
// 16'h665d, 16'h64f9, 16'h6186, 16'h5c19,
// 16'h54d0, 16'h4bce, 16'h4142, 16'h3567,
// 16'h2870, 16'h1ab0, 16'h0c5e, 16'hfdcf,
// 16'hef4e, 16'he11c, 16'hd395, 16'hc6e9,
// 16'hbb70, 16'hb150, 16'ha8d2, 16'ha212,
// 16'h9d3b, 16'h9a65, 16'h999e, 16'h9ae9,
// 16'h9e44, 16'ha392, 16'haacb, 16'hb3b2,
// 16'hbe31, 16'hc9f9, 16'hd6e5, 16'he49b,
// 16'hf2ea, 16'h0174, 16'h0ffd, 16'h1e2e,
// 16'h2bc6, 16'h3878, 16'h4409, 16'h4e34,
// 16'h56ce, 16'h5da3, 16'h6292, 16'h6583,
// 16'h6666, 16'h6531, 16'h61f9, 16'h5cb8,
// 16'h559f, 16'h4cc8, 16'h425f, 16'h36a5,
// 16'h29c6, 16'h1c18, 16'h0dcf, 16'hff47,
// 16'hf0bb, 16'he286, 16'hd4e1, 16'hc827,
// 16'hbc80, 16'hb247, 16'ha995, 16'ha2a9,
// 16'h9da2, 16'h9a95, 16'h999a, 16'h9ab1,
// 16'h9dd5, 16'ha2f6, 16'ha9fc, 16'hb2be,
// 16'hbd10, 16'hc8c3, 16'hd58a, 16'he339,
// 16'hf175, 16'hffff, 16'h0e8d, 16'h1cc6,
// 16'h2a75, 16'h373e, 16'h42f1, 16'h4d40,
// 16'h5606, 16'h5d09, 16'h622a, 16'h6551,
// 16'h6665, 16'h656b, 16'h625f, 16'h5d56,
// 16'h566b, 16'h4dba, 16'h437e, 16'h37db,
// 16'h2b1d, 16'h1d7d, 16'h0f42, 16'h20bb,
// 16'hf22f, 16'he3ea, 16'hd638, 16'hc95d,
// 16'hbda0, 16'hb337, 16'haa65, 16'ha341,
// 16'h9e0e, 16'h9acb, 16'h999b, 16'h9a7f,
// 16'h9d6a, 16'ha260, 16'ha931, 16'hb1cc,
// 16'hbbf8, 16'hc786, 16'hd43d, 16'he1cd,
// 16'hf00a, 16'hfe85, 16'h0d1c, 16'h1b60,
// 16'h291f, 16'h3602, 16'h41d6, 16'h4c47,
// 16'h553a, 16'h5c6b, 16'h61bb, 16'h651c,
// 16'h665c, 16'h65a0, 16'h62c1, 16'h5def,
// 16'h5730, 16'h4ead, 16'h4493, 16'h3914,
// 16'h2c6e, 16'h1ee1, 16'h10b4, 16'h0230,
// 16'hf3a3, 16'he54f, 16'hd791, 16'hca98,
// 16'hbebe, 16'hb434, 16'hab2d, 16'ha3e9,
// 16'h9e79, 16'h9b08, 16'h99a3, 16'h9a4c,
// 16'h9d0d, 16'ha1c7, 16'ha870, 16'hb0db,
// 16'hbae3, 16'hc651, 16'hd2ea, 16'he06d,
// 16'hee95, 16'hfd12, 16'h0baa, 16'h19f4,
// 16'h27cc, 16'h34c2, 16'h40b3, 16'h4b51,
// 16'h5464, 16'h5bcc, 16'h6147, 16'h64dd,
// 16'h6654, 16'h65cc, 16'h6320, 16'h5e83,
// 16'h57ef, 16'h4f9d, 16'h45a4, 16'h3a4b,
// 16'h2dbb, 16'h2046, 16'h1223, 16'h03a6,
// 16'hf514, 16'he6bc, 16'hd8e5, 16'hcbdc,
// 16'hbfdd, 16'hb530, 16'hac04, 16'ha48c,
// 16'h9eee, 16'h9b4a, 16'h99ab, 16'h9a2a,
// 16'h9ca8, 16'ha13e, 16'ha7aa, 16'haff5,
// 16'hb9d0, 16'hc51d, 16'hd19e, 16'hdf07,
// 16'hed28, 16'hfb9e, 16'h0a32, 16'h1891,
// 16'h266b, 16'h3387, 16'h3f8c, 16'h4a54,
// 16'h538f, 16'h5b20, 16'h60d6, 16'h6493,
// 16'h664c, 16'h65ec, 16'h6380, 16'h5f0d,
// 16'h58af, 16'h5083, 16'h46b6, 16'h3b7a,
// 16'h2f0b, 16'h21a6, 16'h1393, 16'h051b,
// 16'hf686, 16'he829, 16'hda3e, 16'hcd1f,
// 16'hc102, 16'hb630, 16'hacdd, 16'ha535,
// 16'h9f6a, 16'h9b8d, 16'h99c0, 16'h9a01,
// 16'h9c55, 16'ha0ae, 16'ha6f5, 16'haf0a,
// 16'hb8c3, 16'hc3ee, 16'hd04f, 16'hddab,
// 16'hebb5, 16'hfa2b, 16'h08bf, 16'h1722,
// 16'h2515, 16'h323e, 16'h3e6a, 16'h494d,
// 16'h52b7, 16'h5a74, 16'h6058, 16'h644d,
// 16'h6635, 16'h6610, 16'h63d4, 16'h5f98,
// 16'h5964, 16'h516a, 16'h47c1, 16'h3caa,
// 16'h3055, 16'h2306, 16'h1501, 16'h0690,
// 16'hf7fa, 16'he995, 16'hdb99, 16'hce66,
// 16'hc229, 16'hb737, 16'hadb6, 16'ha5e7,
// 16'h9fe6, 16'h9bd9, 16'h99d8, 16'h99e1,
// 16'h9c03, 16'ha027, 16'ha63f, 16'hae28,
// 16'hb7b7, 16'hc2c3, 16'hcf04, 16'hdc4e,
// 16'hea46, 16'hf8b6, 16'h074c, 16'h15b5,
// 16'h23b8, 16'h30f7, 16'h3d40, 16'h4847,
// 16'h51da, 16'h59bf, 16'h5fda, 16'h63fe,
// 16'h661b, 16'h662e, 16'h6422, 16'h601c,
// 16'h5a19, 16'h5249, 16'h48cb, 16'h3dd4,
// 16'h319e, 16'h2462, 16'h1670, 16'h0804,
// 16'hf96f, 16'heb01, 16'hdcf8, 16'hcfac,
// 16'hc358, 16'hb83c, 16'hae99, 16'ha69a,
// 16'ha068, 16'h9c2d, 16'h99f0, 16'h99ca,
// 16'h9bb5, 16'h9fa6, 16'ha58e, 16'had47,
// 16'hb6b5, 16'hc194, 16'hcdc3, 16'hdaeb,
// 16'he8de, 16'hf740, 16'h05d6, 16'h144b,
// 16'h2255, 16'h2fb0, 16'h3c13, 16'h473b,
// 16'h50f9, 16'h5908, 16'h5f56, 16'h63a7,
// 16'h6602, 16'h663e, 16'h6473, 16'h6097,
// 16'h5aca, 16'h5324, 16'h49d1, 16'h3efb,
// 16'h32e3, 16'h25c0, 16'h17d9, 16'h097a,
// 16'hfae5, 16'hec6b, 16'hde5d, 16'hd0f2,
// 16'hc488, 16'hb949, 16'haf7d, 16'ha752,
// 16'ha0f3, 16'h9c7e, 16'h9a16, 16'h99b2,
// 16'h9b6f, 16'h9f29, 16'ha4e0, 16'hac71,
// 16'hb5ad, 16'hc072, 16'hcc7b, 16'hd993,
// 16'he771, 16'hf5ce, 16'h0460, 16'h12db,
// 16'h20f5, 16'h2e65, 16'h3ae3, 16'h462e,
// 16'h500f, 16'h5850, 16'h5ec7, 16'h6355,
// 16'h65d8, 16'h6655, 16'h64b4, 16'h6115,
// 16'h5b70, 16'h5420, 16'h4ace, 16'h4024,
// 16'h3422, 16'h271d, 16'h1942, 16'h0aef,
// 16'hfc57, 16'heddf, 16'hdfb9, 16'hd245,
// 16'hc5b6, 16'hba59, 16'hb067, 16'ha80e,
// 16'ha17f, 16'h9cde, 16'h9a36, 16'h99aa,
// 16'h9b26, 16'h9eb4, 16'ha438, 16'hab9b,
// 16'hb4ae, 16'hbf50, 16'hcb38, 16'hd83b,
// 16'he607, 16'hf459, 16'h02ed, 16'h116a,
// 16'h1f94, 16'h2d16, 16'h39af, 16'h451d,
// 16'h4f24, 16'h5791, 16'h5e38, 16'h62f5,
// 16'h65b2, 16'h665d, 16'h64f9, 16'h6185,
// 16'h5c1b, 16'h54ce, 16'h4bcf, 16'h4144,
// 16'h3561, 16'h2879, 16'h1aa7, 16'h0c63,
// 16'hfdcf, 16'hef4a, 16'he123, 16'hd38e,
// 16'hc6ef, 16'hbb6a, 16'hb156, 16'ha8cd,
// 16'ha216, 16'h9d37, 16'h9a6a, 16'h9999,
// 16'h9aee, 16'h9e3e, 16'ha398, 16'haac7,
// 16'hb3b4, 16'hbe30, 16'hc9f9, 16'hd6e5,
// 16'he49c, 16'hf2e9, 16'h0175, 16'h0ffc,
// 16'h1e2d, 16'h2bc8, 16'h3877, 16'h440a,
// 16'h4e33, 16'h56ce, 16'h5da3, 16'h6292,
// 16'h6584, 16'h6664, 16'h6534, 16'h61f6,
// 16'h5cb9, 16'h55a0, 16'h4cc7, 16'h4260,
// 16'h36a4, 16'h29c7, 16'h1c17, 16'h0dd0,
// 16'hff47, 16'hf0bb, 16'he286, 16'hd4e2,
// 16'hc824, 16'hbc84, 16'hb244, 16'ha997,
// 16'ha2a9, 16'h9da1, 16'h9a96, 16'h9999,
// 16'h9ab2, 16'h9dd5, 16'ha2f6, 16'ha9fc,
// 16'hb2bd, 16'hbd12, 16'hc8c1, 16'hd58b,
// 16'he338, 16'hf177, 16'hfffd, 16'h0e8e,
// 16'h1cc5, 16'h2a76, 16'h373e, 16'h42f1,
// 16'h4d3f, 16'h5608, 16'h5d06, 16'h622d,
// 16'h654f, 16'h6665, 16'h656c, 16'h625e,
// 16'h5d56, 16'h566b, 16'h4dbb, 16'h437c,
// 16'h37de, 16'h2b1a, 16'h1d7f, 16'h0f41,
// 16'h20bc, 16'hf22e, 16'he3ea, 16'hd638,
// 16'hc95e, 16'hbd9e, 16'hb33a, 16'haa60,
// 16'ha346, 16'h9e0b, 16'h9acc, 16'h999b,
// 16'h9a7e, 16'h9d6b, 16'ha260, 16'ha931,
// 16'hb1cb, 16'hbbf9, 16'hc786, 16'hd43b,
// 16'he1d2, 16'hf003, 16'hfe8b, 16'h0d18,
// 16'h1b63, 16'h291d, 16'h3604, 16'h41d3,
// 16'h4c49, 16'h553b, 16'h5c68, 16'h61c0,
// 16'h6516, 16'h6661, 16'h659d, 16'h62c3,
// 16'h5dee, 16'h5731, 16'h4eab, 16'h4495,
// 16'h3913, 16'h2c6f, 16'h1ee0, 16'h10b5,
// 16'h022f, 16'hf3a2, 16'he552, 16'hd78d,
// 16'hca9c, 16'hbebc, 16'hb433, 16'hab2f,
// 16'ha3e7, 16'h9e7a, 16'h9b09, 16'h99a1,
// 16'h9a4e, 16'h9d0c, 16'ha1c7, 16'ha870,
// 16'hb0dc, 16'hbae2, 16'hc652, 16'hd2e9,
// 16'he06d, 16'hee95, 16'hfd14, 16'h0ba6,
// 16'h19f9, 16'h27c7, 16'h34c5, 16'h40b4,
// 16'h4b4e, 16'h5467, 16'h5bc9, 16'h6149,
// 16'h64dd, 16'h6654, 16'h65cb, 16'h6321,
// 16'h5e83, 16'h57ef, 16'h4f9c, 16'h45a5,
// 16'h3a4a, 16'h2dbe, 16'h2042, 16'h1227,
// 16'h03a2, 16'hf518, 16'he6b8, 16'hd8e8,
// 16'hcbda, 16'hbfdf, 16'hb530, 16'hac01,
// 16'ha48f, 16'h9eec, 16'h9b4c, 16'h99ab,
// 16'h9a27, 16'h9cad, 16'ha138, 16'ha7b1,
// 16'hafef, 16'hb9d2, 16'hc51f, 16'hd19a,
// 16'hdf0c, 16'hed24, 16'hfb9f, 16'h0a34,
// 16'h188e, 16'h266e, 16'h3384, 16'h3f90,
// 16'h4a50, 16'h5392, 16'h5b1f, 16'h60d5,
// 16'h6496, 16'h6648, 16'h65f0, 16'h637c,
// 16'h5f11, 16'h58ab, 16'h5086, 16'h46b4,
// 16'h3b7d, 16'h2f07, 16'h21a9, 16'h1391,
// 16'h051c, 16'hf688, 16'he824, 16'hda42,
// 16'hcd1c, 16'hc105, 16'hb630, 16'hacda,
// 16'ha537, 16'h9f69, 16'h9b8e, 16'h99c0,
// 16'h9a01, 16'h9c54, 16'ha0b0, 16'ha6f3,
// 16'haf0b, 16'hb8c3, 16'hc3ed, 16'hd051,
// 16'hdda9, 16'hebb7, 16'hfa29, 16'h08c0,
// 16'h1723, 16'h2512, 16'h3242, 16'h3e66,
// 16'h4950, 16'h52b6, 16'h5a73, 16'h6059,
// 16'h644c, 16'h6636, 16'h660f, 16'h63d5,
// 16'h5f96, 16'h5966, 16'h5169, 16'h47c1,
// 16'h3caa, 16'h3055, 16'h2306, 16'h1501,
// 16'h068f, 16'hf7fc, 16'he992, 16'hdb9d,
// 16'hce63, 16'hc22a, 16'hb736, 16'hadb8,
// 16'ha5e5, 16'h9fe7, 16'h9bda, 16'h99d5,
// 16'h99e5, 16'h9c20, 16'ha029, 16'ha63d,
// 16'hae29, 16'hb7b8, 16'hc2c1, 16'hcf08,
// 16'hdc49, 16'hea4a, 16'hf8b4, 16'h074c,
// 16'h15b5, 16'h23b9, 16'h30f5, 16'h3d43,
// 16'h4844, 16'h51db, 16'h59c0, 16'h5fd8,
// 16'h63ff, 16'h661c, 16'h662b, 16'h6427,
// 16'h6016, 16'h5a1e, 16'h5245, 16'h48ce,
// 16'h3dd2, 16'h319f, 16'h2462, 16'h166f,
// 16'h0805, 16'hf96e, 16'heb01, 16'hdcf9,
// 16'hcfac, 16'hc356, 16'hb83f, 16'hae96,
// 16'ha69c, 16'ha067, 16'h9c2d, 16'h99f1,
// 16'h99c9, 16'h9bb5, 16'h9fa6, 16'ha58e,
// 16'had49, 16'hb6b2, 16'hc196, 16'hcdc2,
// 16'hdaed, 16'he8db, 16'hf744, 16'h05d2,
// 16'h144e, 16'h2253, 16'h2fb2, 16'h3c11,
// 16'h473d, 16'h50f6, 16'h590c, 16'h5f51,
// 16'h63ad, 16'h65fb, 16'h6644, 16'h646f,
// 16'h6099, 16'h5aca, 16'h5323, 16'h49d1,
// 16'h3efb, 16'h32e5, 16'h25bd, 16'h17dd,
// 16'h0975, 16'hfae8, 16'hec6b, 16'hde5b,
// 16'hd0f5, 16'hc486, 16'hb94a, 16'haf7c,
// 16'ha752, 16'ha0f2, 16'h9c81, 16'h9a13,
// 16'h99b5, 16'h9b6c, 16'h9f2a, 16'ha4e1,
// 16'hac6f, 16'hb5ae, 16'hc072, 16'hcc7b,
// 16'hd994, 16'he76e, 16'hf5d0, 16'h045e,
// 16'h12de, 16'h20f4, 16'h2e65, 16'h3ae0,
// 16'h4632, 16'h500c, 16'h5854, 16'h5ec4,
// 16'h6355, 16'h65d9, 16'h6654, 16'h64b6,
// 16'h6111, 16'h5b75, 16'h53fc, 16'h4ad0,
// 16'h4023, 16'h3424, 16'h271a, 16'h1946,
// 16'h0aea, 16'hfc5b, 16'hedde, 16'hdfb9,
// 16'hd244, 16'hc5b7, 16'hba59, 16'hb066,
// 16'ha810, 16'ha17e, 16'h9cdc, 16'h9a3a,
// 16'h99a7, 16'h9b27, 16'h9eb6, 16'ha435,
// 16'hab9c, 16'hb4b0, 16'hbf4c, 16'hcb3d,
// 16'hd837, 16'he607, 16'hf45c, 16'h02e9,
// 16'h116e, 16'h1f91, 16'h2d18, 16'h39ad,
// 16'h451e, 16'h4f25, 16'h578f, 16'h5e3b,
// 16'h62f1, 16'h65b5, 16'h665b, 16'h64fb,
// 16'h6183, 16'h5c1c, 16'h54ce, 16'h4bcf,
// 16'h4143, 16'h3563, 16'h2876, 16'h1aaa,
// 16'h0c63, 16'hfdcb, 16'hef51, 16'he11a,
// 16'hd397, 16'hc6e8, 16'hbb6f, 16'hb152,
// 16'ha8d0, 16'ha214, 16'h9d3a, 16'h9a66,
// 16'h999d, 16'h9aea, 16'h9e42, 16'ha396,
// 16'haac7, 16'hb3b6, 16'hbe2d, 16'hc9fc,
// 16'hd6e2, 16'he49f, 16'hf2e7, 16'h0176,
// 16'h0ffc, 16'h1e2d, 16'h2bc8, 16'h3877,
// 16'h4409, 16'h4e34, 16'h56ce, 16'h5da2,
// 16'h6294, 16'h6582, 16'h6665, 16'h6534,
// 16'h61f4, 16'h5cbc, 16'h559f, 16'h4cc5,
// 16'h4264, 16'h369f, 16'h29cc, 16'h1c13,
// 16'h0dd3, 16'hff43, 16'hf0bf, 16'he283,
// 16'hd4e4, 16'hc823, 16'hbc84, 16'hb243,
// 16'ha999, 16'ha2a6, 16'h9da4, 16'h9a94,
// 16'h999b, 16'h9aaf, 16'h9dd8, 16'ha2f3,
// 16'haa20, 16'hb2b9, 16'hbd15, 16'hc8be,
// 16'hd58f, 16'he335, 16'hf178, 16'hfffd,
// 16'h0e8e, 16'h1cc6, 16'h2a74, 16'h3741,
// 16'h42ed, 16'h4d43, 16'h5605, 16'h5d08,
// 16'h622c, 16'h6550, 16'h6663, 16'h656f,
// 16'h625b, 16'h5d59, 16'h5669, 16'h4dba,
// 16'h437f, 16'h37db, 16'h2b1d, 16'h1d7c,
// 16'h0f42, 16'h20bc, 16'hf22e, 16'he3eb,
// 16'hd636, 16'hc960, 16'hbd9c, 16'hb33c,
// 16'haa5e, 16'ha349, 16'h9e07, 16'h9ad0,
// 16'h9998, 16'h9a7f, 16'h9d6d, 16'ha25c,
// 16'ha935, 16'hb1c8, 16'hbbfb, 16'hc785,
// 16'hd43c, 16'he1d0, 16'hf005, 16'hfe8a,
// 16'h0d1a, 16'h1b60, 16'h291f, 16'h3603,
// 16'h41d3, 16'h4c4b, 16'h5538, 16'h5c6a,
// 16'h61bf, 16'h6516, 16'h6663, 16'h6599,
// 16'h62c7, 16'h5deb, 16'h5732, 16'h4ead,
// 16'h4492, 16'h3915, 16'h2c6e, 16'h1ee0,
// 16'h10b6, 16'h022f, 16'hf3a1, 16'he552,
// 16'hd78e, 16'hca9b, 16'hbebd, 16'hb433,
// 16'hab2e, 16'ha3e8, 16'h9e7a, 16'h9b07,
// 16'h99a4, 16'h9a4c, 16'h9d0d, 16'ha1c7,
// 16'ha86f, 16'hb0dd, 16'hbae1, 16'hc654,
// 16'hd2e6, 16'he071, 16'hee91, 16'hfd16,
// 16'h0ba7, 16'h19f6, 16'h27cb, 16'h34c2,
// 16'h40b4, 16'h4b50, 16'h5466, 16'h5bc9,
// 16'h614a, 16'h64da, 16'h6658, 16'h65c8,
// 16'h6323, 16'h5e81, 16'h57f0, 16'h4f9d,
// 16'h45a3, 16'h3a4c, 16'h2dba, 16'h2047,
// 16'h1223, 16'h03a6, 16'hf513, 16'he6bd,
// 16'hd8e4, 16'hcbdc, 16'hbfe0, 16'hb52b,
// 16'hac09, 16'ha487, 16'h9ef3, 16'h9b46,
// 16'h99af, 16'h9a25, 16'h9cad, 16'ha13a,
// 16'ha7ae, 16'haff2, 16'hb9d0, 16'hc520,
// 16'hd199, 16'hdf0d, 16'hed22, 16'hfba2,
// 16'h0a31, 16'h1890, 16'h266d, 16'h3384,
// 16'h3f8f, 16'h4a52, 16'h5390, 16'h5b20,
// 16'h60d5, 16'h6495, 16'h6649, 16'h65f0,
// 16'h637d, 16'h5f0e, 16'h58af, 16'h5082,
// 16'h46b8, 16'h3b79, 16'h2f0b, 16'h21a5,
// 16'h1395, 16'h0519, 16'hf689, 16'he826,
// 16'hda3f, 16'hcd1f, 16'hc102, 16'hb631,
// 16'hacdc, 16'ha536, 16'h9f68, 16'h9b8e,
// 16'h99c0, 16'h9a01, 16'h9c56, 16'ha0ad,
// 16'ha6f5, 16'haf09, 16'hb8c4, 16'hc3ed,
// 16'hd052, 16'hdda8, 16'hebb6, 16'hfa2c,
// 16'h08bb, 16'h1729, 16'h250d, 16'h3245,
// 16'h3e65, 16'h4950, 16'h52b6, 16'h5a73,
// 16'h605a, 16'h644b, 16'h6637, 16'h660f,
// 16'h63d4, 16'h5f98, 16'h5963, 16'h516c,
// 16'h47bf, 16'h3cac, 16'h3053, 16'h2307,
// 16'h1520, 16'h0691, 16'hf7fa, 16'he994,
// 16'hdb9b, 16'hce63, 16'hc22c, 16'hb734,
// 16'hadb9, 16'ha5e5, 16'h9fe6, 16'h9bdb,
// 16'h99d5, 16'h99e2, 16'h9c04, 16'ha026,
// 16'ha640, 16'hae27, 16'hb7b7, 16'hc2c3,
// 16'hcf06, 16'hdc4a, 16'hea4b, 16'hf8b2,
// 16'h074e, 16'h15b5, 16'h23b6, 16'h30fa,
// 16'h3d3e, 16'h4849, 16'h51d6, 16'h59c3,
// 16'h5fd8, 16'h63fe, 16'h661e, 16'h6628,
// 16'h6428, 16'h6018, 16'h5a1c, 16'h5247,
// 16'h48cb, 16'h3dd6, 16'h319a, 16'h2468,
// 16'h166a, 16'h0807, 16'hf96f, 16'heaff,
// 16'hdcfb, 16'hcfaa, 16'hc358, 16'hb83d,
// 16'hae98, 16'ha69a, 16'ha06a, 16'h9c2a,
// 16'h99f3, 16'h99c7, 16'h9bb8, 16'h9fa3,
// 16'ha591, 16'had45, 16'hb6b6, 16'hc193,
// 16'hcdc4, 16'hdaeb, 16'he8de, 16'hf740,
// 16'h05d6, 16'h144a, 16'h2257, 16'h2faf,
// 16'h3c13, 16'h473c, 16'h50f7, 16'h590b,
// 16'h5f52, 16'h63ab, 16'h65fe, 16'h6642,
// 16'h6470, 16'h6098, 16'h5aca, 16'h5324,
// 16'h49d0, 16'h3efd, 16'h32e1, 16'h25c2,
// 16'h17d8, 16'h097a, 16'hfae4, 16'hec6e,
// 16'hde5a, 16'hd0f5, 16'hc486, 16'hb949,
// 16'haf7e, 16'ha750, 16'ha0f5, 16'h9c7e,
// 16'h9a14, 16'h99b6, 16'h9b69, 16'h9f2e,
// 16'ha4dd, 16'hac73, 16'hb5ab, 16'hc075,
// 16'hcc78, 16'hd995, 16'he770, 16'hf5ce,
// 16'h0460, 16'h12dc, 16'h20f4, 16'h2e66,
// 16'h3ae2, 16'h462d, 16'h5011, 16'h584f,
// 16'h5ec8, 16'h6354, 16'h65d8, 16'h6655,
// 16'h64b5, 16'h6113, 16'h5b73, 16'h53fd,
// 16'h4ad0, 16'h4022, 16'h3425, 16'h271a,
// 16'h1945, 16'h0aeb, 16'hfc5a, 16'hedde,
// 16'hdfba, 16'hd244, 16'hc5b6, 16'hba5a,
// 16'hb065, 16'ha811, 16'ha17d, 16'h9cde,
// 16'h9a38, 16'h99a6, 16'h9b2a, 16'h9eb2,
// 16'ha439, 16'hab9a, 16'hb4b0, 16'hbf4c,
// 16'hcb3d, 16'hd837, 16'he609, 16'hf459,
// 16'h02eb, 16'h116c, 16'h1f94, 16'h2d14,
// 16'h39b2, 16'h4519, 16'h4f28, 16'h578f,
// 16'h5e38, 16'h62f5, 16'h65b2, 16'h665e,
// 16'h64f8, 16'h6186, 16'h5c19, 16'h54d0,
// 16'h4bcf, 16'h4142, 16'h3565, 16'h2873,
// 16'h1aac, 16'h0c61, 16'hfdcf, 16'hef4c,
// 16'he11f, 16'hd393, 16'hc6e8, 16'hbb73,
// 16'hb14c, 16'ha8d6, 16'ha20f, 16'h9d3d,
// 16'h9a65, 16'h999d, 16'h9aea, 16'h9e42,
// 16'ha395, 16'haaca, 16'hb3b2, 16'hbe31,
// 16'hc9f9, 16'hd6e4, 16'he49e, 16'hf2e7,
// 16'h0177, 16'h0ff9, 16'h1e32, 16'h2bc2,
// 16'h387d, 16'h4404, 16'h4e38, 16'h56cb,
// 16'h5da4, 16'h6292, 16'h6584, 16'h6664,
// 16'h6534, 16'h61f5, 16'h5cba, 16'h55a0,
// 16'h4cc6, 16'h4262, 16'h36a1, 16'h29ca,
// 16'h1c14, 16'h0dd3, 16'hff44, 16'hf0be,
// 16'he283, 16'hd4e4, 16'hc823, 16'hbc84,
// 16'hb245, 16'ha995, 16'ha2ac, 16'h9d9d,
// 16'h9a99, 16'h9998, 16'h9ab1, 16'h9dd7,
// 16'ha2f4, 16'ha9fe, 16'hb2bb, 16'hbd14,
// 16'hc8be, 16'hd58e, 16'he338, 16'hf174,
// 16'h2002, 16'h0e89, 16'h1cc9, 16'h2a73,
// 16'h3741, 16'h42ed, 16'h4d44, 16'h5604,
// 16'h5d08, 16'h622e, 16'h654b, 16'h666a,
// 16'h6568, 16'h6260, 16'h5d56, 16'h566a,
// 16'h4dbc, 16'h437c, 16'h37dd, 16'h2b1b,
// 16'h1d7e, 16'h0f42, 16'h20bb, 16'hf22f,
// 16'he3ea, 16'hd637, 16'hc95f, 16'hbd9c,
// 16'hb33d, 16'haa5d, 16'ha349, 16'h9e09,
// 16'h9acc, 16'h999c, 16'h9a7c, 16'h9d6f,
// 16'ha25c, 16'ha934, 16'hb1c9, 16'hbbfa,
// 16'hc785, 16'hd43e, 16'he1cd, 16'hf009,
// 16'hfe86, 16'h0d1b, 16'h1b61, 16'h291e,
// 16'h3604, 16'h41d3, 16'h4c49, 16'h553b,
// 16'h5c68, 16'h61c0, 16'h6515, 16'h6663,
// 16'h659b, 16'h62c4, 16'h5def, 16'h572e,
// 16'h4eae, 16'h4494, 16'h3912, 16'h2c71,
// 16'h1ede, 16'h10b7, 16'h022d, 16'hf3a5,
// 16'he54d, 16'hd793, 16'hca96, 16'hbec1,
// 16'hb430, 16'hab31, 16'ha3e6, 16'h9e7a,
// 16'h9b08, 16'h99a3, 16'h9a4d, 16'h9d0c,
// 16'ha1c8, 16'ha86e, 16'hb0de, 16'hbae0,
// 16'hc653, 16'hd2ea, 16'he06b, 16'hee98,
// 16'hfd10, 16'h0baa, 16'h19f6, 16'h27c9,
// 16'h34c4, 16'h40b3, 16'h4b51, 16'h5464,
// 16'h5bca, 16'h614a, 16'h64db, 16'h6656,
// 16'h65c9, 16'h6322, 16'h5e83, 16'h57ef,
// 16'h4f9c, 16'h45a5, 16'h3a49, 16'h2dbe,
// 16'h2044, 16'h1224, 16'h03a6, 16'hf514,
// 16'he6ba, 16'hd8e8, 16'hcbd9, 16'hbfe0,
// 16'hb52e, 16'hac05, 16'ha48a, 16'h9ef1,
// 16'h9b47, 16'h99af, 16'h9a25, 16'h9cad,
// 16'ha13a, 16'ha7ae, 16'haff2, 16'hb9d1,
// 16'hc51e, 16'hd19c, 16'hdf0a, 16'hed25,
// 16'hfb9f, 16'h0a34, 16'h188d, 16'h2670,
// 16'h3382, 16'h3f90, 16'h4a51, 16'h5390,
// 16'h5b22, 16'h60d2, 16'h6498, 16'h6647,
// 16'h65f0, 16'h637e, 16'h5f0e, 16'h58ae,
// 16'h5084, 16'h46b5, 16'h3b7c, 16'h2f09,
// 16'h21a7, 16'h1393, 16'h051a, 16'hf688,
// 16'he826, 16'hda40, 16'hcd1e, 16'hc103,
// 16'hb630, 16'hacdc, 16'ha536, 16'h9f68,
// 16'h9b8f, 16'h99bf, 16'h9a02, 16'h9c54,
// 16'ha0af, 16'ha6f3, 16'haf0c, 16'hb8c2,
// 16'hc3ee, 16'hd051, 16'hdda8, 16'hebb8,
// 16'hfa28, 16'h08c1, 16'h1722, 16'h2514,
// 16'h323e, 16'h3e6b, 16'h494c, 16'h52b8,
// 16'h5a73, 16'h6057, 16'h644f, 16'h6634,
// 16'h6610, 16'h63d4, 16'h5f97, 16'h5966,
// 16'h5168, 16'h47c3, 16'h3ca8, 16'h3057,
// 16'h2303, 16'h1504, 16'h068c, 16'hf820,
// 16'he98f, 16'hdb9e, 16'hce61, 16'hc22d,
// 16'hb734, 16'hadb8, 16'ha5e6, 16'h9fe6,
// 16'h9bdb, 16'h99d5, 16'h99e3, 16'h9c02,
// 16'ha028, 16'ha63e, 16'hae28, 16'hb7b8,
// 16'hc2c2, 16'hcf06, 16'hdc4c, 16'hea46,
// 16'hf8b8, 16'h0749, 16'h15b8, 16'h23b6,
// 16'h30f7, 16'h3d42, 16'h4845, 16'h51da,
// 16'h59c0, 16'h5fd9, 16'h63fe, 16'h661d,
// 16'h662a, 16'h6425, 16'h601b, 16'h5a19,
// 16'h524a, 16'h48ca, 16'h3dd4, 16'h319e,
// 16'h2462, 16'h1672, 16'h0820, 16'hf974,
// 16'heafc, 16'hdcfc, 16'hcfaa, 16'hc358,
// 16'hb83d, 16'hae98, 16'ha69a, 16'ha069,
// 16'h9c2b, 16'h99f3, 16'h99c8, 16'h9bb5,
// 16'h9fa6, 16'ha58e, 16'had49, 16'hb6b2,
// 16'hc198, 16'hcdbe, 16'hdaf0, 16'he8da,
// 16'hf743, 16'h05d5, 16'h144a, 16'h2256,
// 16'h2fb0, 16'h3c12, 16'h473e, 16'h50f4,
// 16'h590d, 16'h5f51, 16'h63ac, 16'h65fe,
// 16'h6641, 16'h6471, 16'h6098, 16'h5aca,
// 16'h5323, 16'h49d2, 16'h3efa, 16'h32e5,
// 16'h25bd, 16'h17dd, 16'h0976, 16'hfae6,
// 16'hec6d, 16'hde59, 16'hd0f8, 16'hc482,
// 16'hb94d, 16'haf7a, 16'ha754, 16'ha0f1,
// 16'h9c81, 16'h9a13, 16'h99b5, 16'h9b6d,
// 16'h9f29, 16'ha4e1, 16'hac70, 16'hb5ae,
// 16'hc072, 16'hcc7b, 16'hd993, 16'he770,
// 16'hf5cf, 16'h045f, 16'h12dd, 16'h20f4,
// 16'h2e65, 16'h3ae1, 16'h4630, 16'h500f,
// 16'h5850, 16'h5ec8, 16'h6351, 16'h65dd,
// 16'h6650, 16'h64b9, 16'h6110, 16'h5b75,
// 16'h53fb, 16'h4ad3, 16'h401e, 16'h3429,
// 16'h2717, 16'h1946, 16'h0aeb, 16'hfc5c,
// 16'hedda, 16'hdfbd, 16'hd243, 16'hc5b6,
// 16'hba5a, 16'hb066, 16'ha80e, 16'ha181,
// 16'h9cdb, 16'h9a3a, 16'h99a5, 16'h9b2b,
// 16'h9eb1, 16'ha43a, 16'hab99, 16'hb4b0,
// 16'hbf4d, 16'hcb3c, 16'hd838, 16'he608,
// 16'hf459, 16'h02eb, 16'h116d, 16'h1f92,
// 16'h2d17, 16'h39ae, 16'h451e, 16'h4f23,
// 16'h5792, 16'h5e37, 16'h62f5, 16'h65b2,
// 16'h665e, 16'h64f8, 16'h6185, 16'h5c1b,
// 16'h54ce, 16'h4bcf, 16'h4143, 16'h3565,
// 16'h2872, 16'h1aae, 16'h0c5f, 16'hfdd0,
// 16'hef4c, 16'he11f, 16'hd391, 16'hc6ee,
// 16'hbb6a, 16'hb157, 16'ha8cc, 16'ha216,
// 16'h9d39, 16'h9a66, 16'h999e, 16'h9aea,
// 16'h9e40, 16'ha399, 16'haac3, 16'hb3ba,
// 16'hbe2a, 16'hc9fd, 16'hd6e4, 16'he49a,
// 16'hf2ec, 16'h0172, 16'h0ffe, 16'h1e2d,
// 16'h2bc6, 16'h387a, 16'h4406, 16'h4e37,
// 16'h56cb, 16'h5da5, 16'h6291, 16'h6585,
// 16'h6663, 16'h6535, 16'h61f3, 16'h5cbd,
// 16'h559d, 16'h4cc9, 16'h425f, 16'h36a4,
// 16'h29c7, 16'h1c16, 16'h0dd3, 16'hff42,
// 16'hf0c1, 16'he280, 16'hd4e6, 16'hc822,
// 16'hbc86, 16'hb242, 16'ha997, 16'ha2aa,
// 16'h9da0, 16'h9a97, 16'h9999, 16'h9ab1,
// 16'h9dd5, 16'ha2f8, 16'ha9f9, 16'hb2bf,
// 16'hbd12, 16'hc8bf, 16'hd58e, 16'he337,
// 16'hf174, 16'h2003, 16'h0e87, 16'h1ccc,
// 16'h2a70, 16'h3742, 16'h42ee, 16'h4d42,
// 16'h5605, 16'h5d09, 16'h622b, 16'h654f,
// 16'h6666, 16'h656a, 16'h6260, 16'h5d56,
// 16'h566b, 16'h4db9, 16'h437f, 16'h37da,
// 16'h2b1e, 16'h1d7c, 16'h0f43, 16'h20bb,
// 16'hf22f, 16'he3e9, 16'hd638, 16'hc95e,
// 16'hbd9f, 16'hb339, 16'haa61, 16'ha344,
// 16'h9e0e, 16'h9ac9, 16'h999e, 16'h9a7a,
// 16'h9d70, 16'ha25b, 16'ha935, 16'hb1c9,
// 16'hbbf9, 16'hc787, 16'hd43a, 16'he1d3,
// 16'hf002, 16'hfe8d, 16'h0d16, 16'h1b63,
// 16'h291e, 16'h3603, 16'h41d5, 16'h4c47,
// 16'h553b, 16'h5c69, 16'h61bf, 16'h6517,
// 16'h6660, 16'h659d, 16'h62c3, 16'h5df0,
// 16'h572e, 16'h4ead, 16'h4494, 16'h3913,
// 16'h2c6f, 16'h1ee1, 16'h10b3, 16'h0232,
// 16'hf39f, 16'he553, 16'hd78f, 16'hca99,
// 16'hbebf, 16'hb430, 16'hab31, 16'ha3e7,
// 16'h9e7a, 16'h9b07, 16'h99a4, 16'h9a4b,
// 16'h9d0f, 16'ha1c5, 16'ha870, 16'hb0dd,
// 16'hbae1, 16'hc653, 16'hd2e9, 16'he06d,
// 16'hee94, 16'hfd15, 16'h0ba6, 16'h19f9,
// 16'h27c7, 16'h34c5, 16'h40b3, 16'h4b4f,
// 16'h5468, 16'h5bc6, 16'h614d, 16'h64d8,
// 16'h6659, 16'h65c7, 16'h6324, 16'h5e81,
// 16'h57ef, 16'h4f9d, 16'h45a5, 16'h3a49,
// 16'h2dbe, 16'h2043, 16'h1226, 16'h03a3,
// 16'hf517, 16'he6b8, 16'hd8e8, 16'hcbdb,
// 16'hbfdd, 16'hb532, 16'hac20, 16'ha48f,
// 16'h9eec, 16'h9b4c, 16'h99ab, 16'h9a27,
// 16'h9cac, 16'ha13b, 16'ha7ac, 16'haff5,
// 16'hb9cc, 16'hc523, 16'hd198, 16'hdf0e,
// 16'hed21, 16'hfba3, 16'h0a2f, 16'h1893,
// 16'h2669, 16'h3389, 16'h3f8b, 16'h4a55,
// 16'h538e, 16'h5b21, 16'h60d4, 16'h6496,
// 16'h6649, 16'h65ef, 16'h637e, 16'h5f0f,
// 16'h58ac, 16'h5085, 16'h46b5, 16'h3b7c,
// 16'h2f09, 16'h21a7, 16'h1392, 16'h051c,
// 16'hf686, 16'he828, 16'hda3e, 16'hcd1f,
// 16'hc103, 16'hb630, 16'hacdc, 16'ha536,
// 16'h9f68, 16'h9b90, 16'h99be, 16'h9a01,
// 16'h9c58, 16'ha0a8, 16'ha6fc, 16'haf05,
// 16'hb8c4, 16'hc3f0, 16'hd04d, 16'hddac,
// 16'hebb5, 16'hfa2a, 16'h08c0, 16'h1723,
// 16'h2514, 16'h323d, 16'h3e6b, 16'h494c,
// 16'h52ba, 16'h5a70, 16'h605c, 16'h6449,
// 16'h6638, 16'h660e, 16'h63d5, 16'h5f97,
// 16'h5966, 16'h5167, 16'h47c5, 16'h3ca6,
// 16'h3058, 16'h2303, 16'h1503, 16'h068f,
// 16'hf7fc, 16'he992, 16'hdb9c, 16'hce62,
// 16'hc22f, 16'hb730, 16'hadbc, 16'ha5e3,
// 16'h9fe7, 16'h9bdb, 16'h99d5, 16'h99e3,
// 16'h9c03, 16'ha026, 16'ha640, 16'hae27,
// 16'hb7b9, 16'hc2c1, 16'hcf06, 16'hdc4c,
// 16'hea47, 16'hf8b8, 16'h0748, 16'h15b9,
// 16'h23b4, 16'h30fa, 16'h3d3f, 16'h4847,
// 16'h51d9, 16'h59c0, 16'h5fdb, 16'h63fa,
// 16'h6622, 16'h6625, 16'h642a, 16'h6016,
// 16'h5a1e, 16'h5245, 16'h48cf, 16'h3dd0,
// 16'h31a0, 16'h2462, 16'h1670, 16'h0803,
// 16'hf971, 16'heaff, 16'hdcfa, 16'hcfab,
// 16'hc357, 16'hb83d, 16'hae9a, 16'ha698,
// 16'ha06b, 16'h9c29, 16'h99f4, 16'h99c7,
// 16'h9bb7, 16'h9fa4, 16'ha590, 16'had47,
// 16'hb6b3, 16'hc197, 16'hcdc0, 16'hdaee,
// 16'he8dd, 16'hf73f, 16'h05d8, 16'h1448,
// 16'h2258, 16'h2fae, 16'h3c15, 16'h4739,
// 16'h50fa, 16'h5907, 16'h5f56, 16'h63a8,
// 16'h6601, 16'h663f, 16'h6472, 16'h6098,
// 16'h5ac9, 16'h5325, 16'h49d0, 16'h3efc,
// 16'h32e3, 16'h25c0, 16'h17d9, 16'h097b,
// 16'hfae1, 16'hec72, 16'hde54, 16'hd0fc,
// 16'hc480, 16'hb94d, 16'haf7b, 16'ha753,
// 16'ha0f1, 16'h9c82, 16'h9a11, 16'h99b8,
// 16'h9b69, 16'h9f2e, 16'ha4dc, 16'hac73,
// 16'hb5ad, 16'hc072, 16'hcc7c, 16'hd991,
// 16'he772, 16'hf5cc, 16'h0463, 16'h12d8,
// 16'h20f9, 16'h2e61, 16'h3ae5, 16'h462c,
// 16'h5012, 16'h584d, 16'h5ecc, 16'h634e,
// 16'h65de, 16'h6651, 16'h64b7, 16'h6112,
// 16'h5b74, 16'h53fc, 16'h4ad0, 16'h4023,
// 16'h3423, 16'h271d, 16'h1943, 16'h0aeb,
// 16'hfc5c, 16'hedda, 16'hdfbf, 16'hd23f,
// 16'hc5b9, 16'hba5a, 16'hb064, 16'ha810,
// 16'ha180, 16'h9cda, 16'h9a3b, 16'h99a6,
// 16'h9b28, 16'h9eb4, 16'ha438, 16'hab9a,
// 16'hb4af, 16'hbf50, 16'hcb37, 16'hd83c,
// 16'he606, 16'hf45a, 16'h02ed, 16'h1169,
// 16'h1f94, 16'h2d17, 16'h39ae, 16'h451e,
// 16'h4f23, 16'h5792, 16'h5e36, 16'h62f7,
// 16'h65b0, 16'h665f, 16'h64f8, 16'h6185,
// 16'h5c1b, 16'h54ce, 16'h4bd0, 16'h4141,
// 16'h3566, 16'h2872, 16'h1aae, 16'h0c60,
// 16'hfdcf, 16'hef4b, 16'he120, 16'hd392,
// 16'hc6ec, 16'hbb6d, 16'hb151, 16'ha8d3,
// 16'ha210, 16'h9d3e, 16'h9a62, 16'h99a0,
// 16'h9ae9, 16'h9e42, 16'ha395, 16'haac8,
// 16'hb3b5, 16'hbe2f, 16'hc9fa, 16'hd6e4,
// 16'he49c, 16'hf2ea, 16'h0173, 16'h0ffe,
// 16'h1e2d, 16'h2bc6, 16'h387a, 16'h4406,
// 16'h4e36, 16'h56ce, 16'h5da1, 16'h6295,
// 16'h6581, 16'h6666, 16'h6533, 16'h61f6,
// 16'h5cba, 16'h559f, 16'h4cc7, 16'h4261,
// 16'h36a2, 16'h29ca, 16'h1c13, 16'h0dd4,
// 16'hff44, 16'hf0bc, 16'he287, 16'hd4df,
// 16'hc828, 16'hbc80, 16'hb248, 16'ha993,
// 16'ha2ac, 16'h9d9e, 16'h9a98, 16'h9999,
// 16'h9ab1, 16'h9dd6, 16'ha2f4, 16'ha9ff,
// 16'hb2ba, 16'hbd15, 16'hc8bd, 16'hd58f,
// 16'he336, 16'hf176, 16'h2020, 16'h0e8b,
// 16'h1cc8, 16'h2a73, 16'h3740, 16'h42ee,
// 16'h4d44, 16'h5603, 16'h5d0b, 16'h6229,
// 16'h6551, 16'h6664, 16'h656c, 16'h625f,
// 16'h5d56, 16'h566a, 16'h4dbb, 16'h437d,
// 16'h37dc, 16'h2b1d, 16'h1d7b, 16'h0f45,
// 16'h20b8, 16'hf231, 16'he3e9, 16'hd638,
// 16'hc95e, 16'hbd9e, 16'hb339, 16'haa62,
// 16'ha345, 16'h9e0c, 16'h9acb, 16'h999b,
// 16'h9a7f, 16'h9d6b, 16'ha260, 16'ha930,
// 16'hb1cc, 16'hbbfa, 16'hc784, 16'hd43e,
// 16'he1cd, 16'hf008, 16'hfe89, 16'h0d18,
// 16'h1b63, 16'h291c, 16'h3606, 16'h41d1,
// 16'h4c4c, 16'h5537, 16'h5c6b, 16'h61be,
// 16'h6518, 16'h665f, 16'h65a0, 16'h62be,
// 16'h5df4, 16'h572b, 16'h4eb0, 16'h4491,
// 16'h3915, 16'h2c6f, 16'h1edf, 16'h10b7,
// 16'h022b, 16'hf3a6, 16'he54f, 16'hd790,
// 16'hca9a, 16'hbebc, 16'hb434, 16'hab2f,
// 16'ha3e7, 16'h9e7a, 16'h9b07, 16'h99a4,
// 16'h9a4d, 16'h9d0c, 16'ha1c6, 16'ha872,
// 16'hb0d8, 16'hbae8, 16'hc64c, 16'hd2ee,
// 16'he06a, 16'hee96, 16'hfd14, 16'h0ba6,
// 16'h19f9, 16'h27c7, 16'h34c5, 16'h40b3,
// 16'h4b4f, 16'h5468, 16'h5bc5, 16'h6150,
// 16'h64d4, 16'h665d, 16'h65c4, 16'h6325,
// 16'h5e81, 16'h57f1, 16'h4f9a, 16'h45a7,
// 16'h3a48, 16'h2dbe, 16'h2045, 16'h1223,
// 16'h03a6, 16'hf514, 16'he6bb, 16'hd8e7,
// 16'hcbd9, 16'hbfe1, 16'hb52d, 16'hac05,
// 16'ha48c, 16'h9eed, 16'h9b4c, 16'h99a9,
// 16'h9a2a, 16'h9caa, 16'ha13b, 16'ha7af,
// 16'haff0, 16'hb9d2, 16'hc51d, 16'hd19d,
// 16'hdf09, 16'hed26, 16'hfb9f, 16'h0a32,
// 16'h1890, 16'h266d, 16'h3384, 16'h3f8f,
// 16'h4a51, 16'h5391, 16'h5b20, 16'h60d5,
// 16'h6494, 16'h664c, 16'h65eb, 16'h6382,
// 16'h5f0b, 16'h58b0, 16'h5082, 16'h46b8,
// 16'h3b7a, 16'h2f09, 16'h21a8, 16'h1391,
// 16'h051c, 16'hf688, 16'he825, 16'hda41,
// 16'hcd1d, 16'hc104, 16'hb62f, 16'hacdd,
// 16'ha535, 16'h9f6a, 16'h9b8d, 16'h99c1,
// 16'h99ff, 16'h9c57, 16'ha0ad, 16'ha6f5,
// 16'haf0a, 16'hb8c3, 16'hc3ee, 16'hd050,
// 16'hddaa, 16'hebb5, 16'hfa2c, 16'h08bd,
// 16'h1726, 16'h2510, 16'h3242, 16'h3e67,
// 16'h494f, 16'h52b7, 16'h5a72, 16'h6059,
// 16'h644e, 16'h6634, 16'h6610, 16'h63d4,
// 16'h5f96, 16'h5967, 16'h5169, 16'h47c1,
// 16'h3caa, 16'h3054, 16'h2306, 16'h1502,
// 16'h068f, 16'hf7fb, 16'he995, 16'hdb98,
// 16'hce67, 16'hc228, 16'hb737, 16'hadb7,
// 16'ha5e6, 16'h9fe6, 16'h9bda, 16'h99d6,
// 16'h99e3, 16'h9c01, 16'ha029, 16'ha63d,
// 16'hae29, 16'hb7b9, 16'hc2bf, 16'hcf09,
// 16'hdc48, 16'hea4b, 16'hf8b4, 16'h074d,
// 16'h15b4, 16'h23b8, 16'h30f7, 16'h3d40,
// 16'h4848, 16'h51d7, 16'h59c3, 16'h5fd6,
// 16'h6401, 16'h661a, 16'h662d, 16'h6423,
// 16'h601b, 16'h5a1b, 16'h5247, 16'h48cc,
// 16'h3dd4, 16'h319c, 16'h2466, 16'h166b,
// 16'h0808, 16'hf96c, 16'heb03, 16'hdcf7,
// 16'hcfad, 16'hc356, 16'hb83e, 16'hae97,
// 16'ha69b, 16'ha068, 16'h9c2d, 16'h99f0,
// 16'h99ca, 16'h9bb4, 16'h9fa7, 16'ha58c,
// 16'had4b, 16'hb6b0, 16'hc198, 16'hcdc1,
// 16'hdaed, 16'he8db, 16'hf744, 16'h05d1,
// 16'h144f, 16'h2253, 16'h2fb1, 16'h3c13,
// 16'h473b, 16'h50f7, 16'h590b, 16'h5f52,
// 16'h63ac, 16'h65fd, 16'h6643, 16'h646e,
// 16'h609b, 16'h5ac8, 16'h5324, 16'h49d2,
// 16'h3efa, 16'h32e4, 16'h25bf, 16'h17da,
// 16'h0979, 16'hfae5, 16'hec6d, 16'hde59,
// 16'hd0f8, 16'hc482, 16'hb94e, 16'haf79,
// 16'ha755, 16'ha0ef, 16'h9c84, 16'h9a10,
// 16'h99b8, 16'h9b6a, 16'h9f2b, 16'ha4e0,
// 16'hac70, 16'hb5ae, 16'hc071, 16'hcc7d,
// 16'hd991, 16'he772, 16'hf5cd, 16'h045f,
// 16'h12de, 16'h20f3, 16'h2e67, 16'h3adf,
// 16'h4632, 16'h500c, 16'h5853, 16'h5ec6,
// 16'h6352, 16'h65de, 16'h664e, 16'h64bb,
// 16'h610e, 16'h5b77, 16'h53fa, 16'h4ad4,
// 16'h401e, 16'h3427, 16'h271a, 16'h1944,
// 16'h0aee, 16'hfc58, 16'heddd, 16'hdfbc,
// 16'hd242, 16'hc5b7, 16'hba5b, 16'hb063,
// 16'ha813, 16'ha17b, 16'h9cdf, 16'h9a38,
// 16'h99a6, 16'h9b2b, 16'h9eb0, 16'ha43b,
// 16'hab99, 16'hb4af, 16'hbf50, 16'hcb37,
// 16'hd83d, 16'he604, 16'hf45c, 16'h02eb,
// 16'h116a, 16'h1f96, 16'h2d12, 16'h39b3,
// 16'h451a, 16'h4f26, 16'h5790, 16'h5e38,
// 16'h62f4, 16'h65b4, 16'h665b, 16'h64fb,
// 16'h6183, 16'h5c1c, 16'h54ce, 16'h4bcf,
// 16'h4142, 16'h3566, 16'h2872, 16'h1aae,
// 16'h0c5f, 16'hfdcf, 16'hef4e, 16'he11c,
// 16'hd396, 16'hc6e8, 16'hbb70, 16'hb151,
// 16'ha8d1, 16'ha212, 16'h9d3c, 16'h9a64,
// 16'h999f, 16'h9ae8, 16'h9e44, 16'ha394,
// 16'haac8, 16'hb3b6, 16'hbe2b, 16'hca20,
// 16'hd6df, 16'he4a0, 16'hf2e7, 16'h0175,
// 16'h0ffd, 16'h1e2d, 16'h2bc7, 16'h3878,
// 16'h4409, 16'h4e33, 16'h56cf, 16'h5da1,
// 16'h6294, 16'h6582, 16'h6666, 16'h6533,
// 16'h61f4, 16'h5cbd, 16'h559b, 16'h4ccb,
// 16'h425f, 16'h36a2, 16'h29ca, 16'h1c14,
// 16'h0dd3, 16'hff44, 16'hf0be, 16'he282,
// 16'hd4e6, 16'hc822, 16'hbc85, 16'hb244,
// 16'ha995, 16'ha2ab, 16'h9da0, 16'h9a96,
// 16'h999a, 16'h9ab1, 16'h9dd4, 16'ha2f8,
// 16'ha9fa, 16'hb2bf, 16'hbd11, 16'hc8bf,
// 16'hd58f, 16'he335, 16'hf177, 16'h2020,
// 16'h0e89, 16'h1ccb, 16'h2a71, 16'h3742,
// 16'h42ed, 16'h4d43, 16'h5604, 16'h5d0a,
// 16'h622a, 16'h6551, 16'h6665, 16'h656a,
// 16'h6260, 16'h5d55, 16'h566b, 16'h4dbc,
// 16'h437b, 16'h37de, 16'h2b1b, 16'h1d7d,
// 16'h0f43, 16'h20ba, 16'hf230, 16'he3e9,
// 16'hd639, 16'hc95c, 16'hbda1, 16'hb337,
// 16'haa62, 16'ha345, 16'h9e0b, 16'h9acd,
// 16'h999b, 16'h9a7c, 16'h9d6f, 16'ha25a,
// 16'ha937, 16'hb1c7, 16'hbbfc, 16'hc783,
// 16'hd43e, 16'he1ce, 16'hf008, 16'hfe87,
// 16'h0d1b, 16'h1b5f, 16'h2920, 16'h3603,
// 16'h41d2, 16'h4c4c, 16'h5538, 16'h5c69,
// 16'h61c1, 16'h6512, 16'h6667, 16'h6597,
// 16'h62c8, 16'h5deb, 16'h5731, 16'h4ead,
// 16'h4493, 16'h3915, 16'h2c6d, 16'h1ee2,
// 16'h10b2, 16'h0233, 16'hf39f, 16'he554,
// 16'hd78c, 16'hca9b, 16'hbebe, 16'hb431,
// 16'hab32, 16'ha3e3, 16'h9e7e, 16'h9b05,
// 16'h99a4, 16'h9a4d, 16'h9d0b, 16'ha1c9,
// 16'ha86f, 16'hb0db, 16'hbae3, 16'hc652,
// 16'hd2e8, 16'he070, 16'hee91, 16'hfd17,
// 16'h0ba4, 16'h19fb, 16'h27c5, 16'h34c7,
// 16'h40b1, 16'h4b50, 16'h5468, 16'h5bc6,
// 16'h614d, 16'h64d8, 16'h6658, 16'h65c8,
// 16'h6323, 16'h5e82, 16'h57f0, 16'h4f9a,
// 16'h45a8, 16'h3a46, 16'h2dc0, 16'h2044,
// 16'h1222, 16'h03a8, 16'hf513, 16'he6bb,
// 16'hd8e8, 16'hcbd8, 16'hbfe1, 16'hb52e,
// 16'hac03, 16'ha48e, 16'h9eec, 16'h9b4b,
// 16'h99ad, 16'h9a25, 16'h9cae, 16'ha137,
// 16'ha7b2, 16'hafee, 16'hb9d5, 16'hc51b,
// 16'hd19d, 16'hdf0a, 16'hed25, 16'hfba0,
// 16'h0a32, 16'h188f, 16'h266e, 16'h3383,
// 16'h3f91, 16'h4a4f, 16'h5393, 16'h5b1e,
// 16'h60d5, 16'h6496, 16'h6649, 16'h65ee,
// 16'h6380, 16'h5f0c, 16'h58b0, 16'h5081,
// 16'h46b9, 16'h3b79, 16'h2f0a, 16'h21a7,
// 16'h1392, 16'h051b, 16'hf689, 16'he824,
// 16'hda41, 16'hcd1d, 16'hc104, 16'hb630,
// 16'hacdc, 16'ha535, 16'h9f6a, 16'h9b8d,
// 16'h99c1, 16'h9a20, 16'h9c56, 16'ha0ad,
// 16'ha6f6, 16'haf08, 16'hb8c5, 16'hc3ec,
// 16'hd052, 16'hdda9, 16'hebb5, 16'hfa2c,
// 16'h08bd, 16'h1725, 16'h2513, 16'h323e,
// 16'h3e6c, 16'h4949, 16'h52bc, 16'h5a6f,
// 16'h605c, 16'h644a, 16'h6637, 16'h660f,
// 16'h63d4, 16'h5f98, 16'h5964, 16'h516a,
// 16'h47c2, 16'h3ca9, 16'h3055, 16'h2306,
// 16'h1520, 16'h0691, 16'hf7fc, 16'he990,
// 16'hdb9e, 16'hce62, 16'hc22c, 16'hb735,
// 16'hadb7, 16'ha5e6, 16'h9fe7, 16'h9bda,
// 16'h99d5, 16'h99e3, 16'h9c03, 16'ha027,
// 16'ha63f, 16'hae27, 16'hb7b8, 16'hc2c3,
// 16'hcf05, 16'hdc4c, 16'hea47, 16'hf8b7,
// 16'h0749, 16'h15b9, 16'h23b5, 16'h30f8,
// 16'h3d40, 16'h4847, 16'h51d8, 16'h59c3,
// 16'h5fd7, 16'h63fe, 16'h661e, 16'h6629,
// 16'h6428, 16'h6017, 16'h5a1c, 16'h5248,
// 16'h48cb, 16'h3dd5, 16'h319d, 16'h2461,
// 16'h1673, 16'h07ff, 16'hf975, 16'heafc,
// 16'hdcfb, 16'hcfab, 16'hc357, 16'hb83d,
// 16'hae9a, 16'ha697, 16'ha06c, 16'h9c29,
// 16'h99f3, 16'h99c9, 16'h9bb5, 16'h9fa5,
// 16'ha590, 16'had45, 16'hb6b6, 16'hc194,
// 16'hcdc3, 16'hdaec, 16'he8dc, 16'hf742,
// 16'h05d5, 16'h144b, 16'h2255, 16'h2fb1,
// 16'h3c11, 16'h473f, 16'h50f4, 16'h590c,
// 16'h5f52, 16'h63ac, 16'h65fd, 16'h6643,
// 16'h646e, 16'h609b, 16'h5ac7, 16'h5327,
// 16'h49ce, 16'h3efd, 16'h32e3, 16'h25be,
// 16'h17dc, 16'h0977, 16'hfae5, 16'hec6e,
// 16'hde5a, 16'hd0f4, 16'hc488, 16'hb947,
// 16'haf7f, 16'ha751, 16'ha0f3, 16'h9c80,
// 16'h9a12, 16'h99b8, 16'h9b68, 16'h9f2f,
// 16'ha4dd, 16'hac71, 16'hb5ae, 16'hc071,
// 16'hcc7c, 16'hd993, 16'he770, 16'hf5cf,
// 16'h045e, 16'h12de, 16'h20f3, 16'h2e66,
// 16'h3ae2, 16'h462e, 16'h5011, 16'h584e,
// 16'h5ec9, 16'h6352, 16'h65db, 16'h6653,
// 16'h64b6, 16'h6112, 16'h5b74, 16'h53fc,
// 16'h4ad2, 16'h4020, 16'h3425, 16'h271c,
// 16'h1943, 16'h0aee, 16'hfc57, 16'hedde,
// 16'hdfbb, 16'hd243, 16'hc5b8, 16'hba58,
// 16'hb066, 16'ha80e, 16'ha181, 16'h9cdc,
// 16'h9a38, 16'h99a9, 16'h9b25, 16'h9eb5,
// 16'ha43a, 16'hab97, 16'hb4b3, 16'hbf4a,
// 16'hcb3e, 16'hd837, 16'he608, 16'hf45a,
// 16'h02ea, 16'h116f, 16'h1f8f, 16'h2d1a,
// 16'h39ab, 16'h4521, 16'h4f21, 16'h5794,
// 16'h5e35, 16'h62f6, 16'h65b2, 16'h665e,
// 16'h64f8, 16'h6185, 16'h5c1c, 16'h54cc,
// 16'h4bd2, 16'h413f, 16'h3568, 16'h2872,
// 16'h1aac, 16'h0c61, 16'hfdcd, 16'hef50,
// 16'he11b, 16'hd395, 16'hc6e9, 16'hbb6f,
// 16'hb152, 16'ha8d0, 16'ha213, 16'h9d3b,
// 16'h9a66, 16'h999c, 16'h9aeb, 16'h9e40,
// 16'ha398, 16'haac6, 16'hb3b6, 16'hbe2d,
// 16'hc9fc, 16'hd6e2, 16'he49f, 16'hf2e7,
// 16'h0175, 16'h0ffd, 16'h1e2d, 16'h2bc8,
// 16'h3876, 16'h440a, 16'h4e33, 16'h56d0,
// 16'h5da0, 16'h6295, 16'h6581, 16'h6666,
// 16'h6533, 16'h61f6, 16'h5cba, 16'h559f,
// 16'h4cc7, 16'h4260, 16'h36a4, 16'h29c8,
// 16'h1c15, 16'h0dd3, 16'hff43, 16'hf0bf,
// 16'he281, 16'hd4e8, 16'hc81e, 16'hbc8a,
// 16'hb23e, 16'ha99b, 16'ha2a7, 16'h9da2,
// 16'h9a95, 16'h999b, 16'h9aaf, 16'h9dd7,
// 16'ha2f6, 16'ha9fb, 16'hb2bf, 16'hbd10,
// 16'hc8c1, 16'hd58d, 16'he336, 16'hf178,
// 16'hfffd, 16'h0e8d, 16'h1cc7, 16'h2a74,
// 16'h3740, 16'h42ee, 16'h4d43, 16'h5604,
// 16'h5d0a, 16'h622a, 16'h6551, 16'h6664,
// 16'h656c, 16'h625e, 16'h5d57, 16'h566a,
// 16'h4dbb, 16'h437d, 16'h37dc, 16'h2b1d,
// 16'h1d7c, 16'h0f42, 16'h20bc, 16'hf22e,
// 16'he3eb, 16'hd638, 16'hc95c, 16'hbd9f,
// 16'hb33a, 16'haa61, 16'ha345, 16'h9e0c,
// 16'h9ac9, 16'h99a0, 16'h9a79, 16'h9d6f,
// 16'ha25e, 16'ha930, 16'hb1cf, 16'hbbf5,
// 16'hc788, 16'hd43b, 16'he1d0, 16'hf006,
// 16'hfe8a, 16'h0d17, 16'h1b64, 16'h291b,
// 16'h3607, 16'h41cf, 16'h4c4f, 16'h5534,
// 16'h5c6e, 16'h61bc, 16'h6517, 16'h6662,
// 16'h659c, 16'h62c3, 16'h5def, 16'h572f,
// 16'h4ead, 16'h4494, 16'h3913, 16'h2c6f,
// 16'h1ee0, 16'h10b5, 16'h022f, 16'hf3a2,
// 16'he552, 16'hd78d, 16'hca9d, 16'hbeba,
// 16'hb434, 16'hab30, 16'ha3e5, 16'h9e7e,
// 16'h9b03, 16'h99a6, 16'h9a4c, 16'h9d0c,
// 16'ha1c8, 16'ha86f, 16'hb0dc, 16'hbae2,
// 16'hc653, 16'hd2e7, 16'he071, 16'hee8f,
// 16'hfd1a, 16'h0ba1, 16'h19fd, 16'h27c4,
// 16'h34c7, 16'h40b2, 16'h4b50, 16'h5466,
// 16'h5bc8, 16'h614c, 16'h64d9, 16'h6658,
// 16'h65c7, 16'h6325, 16'h5e7f, 16'h57f2,
// 16'h4f9a, 16'h45a6, 16'h3a4a, 16'h2dbc,
// 16'h2045, 16'h1224, 16'h03a5, 16'hf515,
// 16'he6ba, 16'hd8e8, 16'hcbd9, 16'hbfe0,
// 16'hb52f, 16'hac02, 16'ha48e, 16'h9eee,
// 16'h9b48, 16'h99b0, 16'h9a22, 16'h9cb0,
// 16'ha138, 16'ha7af, 16'haff1, 16'hb9d1,
// 16'hc51f, 16'hd19a, 16'hdf0d, 16'hed22,
// 16'hfba2, 16'h0a30, 16'h1891, 16'h266c,
// 16'h3386, 16'h3f8d, 16'h4a53, 16'h538f,
// 16'h5b21, 16'h60d4, 16'h6496, 16'h6649,
// 16'h65ee, 16'h6380, 16'h5f0c, 16'h58b1,
// 16'h5080, 16'h46b9, 16'h3b79, 16'h2f0a,
// 16'h21a8, 16'h1391, 16'h051c, 16'hf687,
// 16'he826, 16'hda3f, 16'hcd20, 16'hc101,
// 16'hb632, 16'hacdb, 16'ha535, 16'h9f6b,
// 16'h9b8c, 16'h99c2, 16'h99ff, 16'h9c56,
// 16'ha0ae, 16'ha6f5, 16'haf09, 16'hb8c5,
// 16'hc3eb, 16'hd053, 16'hdda8, 16'hebb6,
// 16'hfa2c, 16'h08bc, 16'h1727, 16'h250f,
// 16'h3244, 16'h3e64, 16'h4952, 16'h52b4,
// 16'h5a75, 16'h6057, 16'h644f, 16'h6632,
// 16'h6614, 16'h63cf, 16'h5f9b, 16'h5963,
// 16'h516b, 16'h47c1, 16'h3caa, 16'h3052,
// 16'h230a, 16'h14fd, 16'h0694, 16'hf7f8,
// 16'he994, 16'hdb9b, 16'hce64, 16'hc22b,
// 16'hb735, 16'hadb8, 16'ha5e4, 16'h9fe9,
// 16'h9bd8, 16'h99d8, 16'h99e0, 16'h9c04,
// 16'ha027, 16'ha63e, 16'hae2a, 16'hb7b5,
// 16'hc2c4, 16'hcf05, 16'hdc4b, 16'hea4a,
// 16'hf8b3, 16'h074d, 16'h15b5, 16'h23b8,
// 16'h30f6, 16'h3d42, 16'h4844, 16'h51dc,
// 16'h59bf, 16'h5fda, 16'h63fc, 16'h661e,
// 16'h662b, 16'h6424, 16'h601c, 16'h5a18,
// 16'h524a, 16'h48cb, 16'h3dd4, 16'h319d,
// 16'h2463, 16'h1670, 16'h0803, 16'hf971,
// 16'heafe, 16'hdcfb, 16'hcfa9, 16'hc35b,
// 16'hb839, 16'hae9c, 16'ha696, 16'ha06c,
// 16'h9c2a, 16'h99f2, 16'h99ca, 16'h9bb3,
// 16'h9fa7, 16'ha58e, 16'had48, 16'hb6b4,
// 16'hc194, 16'hcdc4, 16'hdaea, 16'he8de,
// 16'hf741, 16'h05d5, 16'h144c, 16'h2254,
// 16'h2fb1, 16'h3c11, 16'h473e, 16'h50f7,
// 16'h5908, 16'h5f56, 16'h63a8, 16'h6601,
// 16'h6640, 16'h6470, 16'h6099, 16'h5ac9,
// 16'h5326, 16'h49cf, 16'h3efc, 16'h32e2,
// 16'h25c1, 16'h17d8, 16'h097c, 16'hfae1,
// 16'hec70, 16'hde59, 16'hd0f5, 16'hc486,
// 16'hb94a, 16'haf7d, 16'ha750, 16'ha0f6,
// 16'h9c7c, 16'h9a17, 16'h99b3, 16'h9b6d,
// 16'h9f2a, 16'ha4e1, 16'hac6e, 16'hb5b1,
// 16'hc06e, 16'hcc80, 16'hd98e, 16'he775,
// 16'hf5cb, 16'h0461, 16'h12db, 16'h20f7,
// 16'h2e62, 16'h3ae5, 16'h462c, 16'h5010,
// 16'h5852, 16'h5ec5, 16'h6355, 16'h65d8,
// 16'h6654, 16'h64b7, 16'h6110, 16'h5b77,
// 16'h53f9, 16'h4ad3, 16'h4021, 16'h3424,
// 16'h271b, 16'h1945, 16'h0aeb, 16'hfc5c,
// 16'hedda, 16'hdfbe, 16'hd23f, 16'hc5bb,
// 16'hba57, 16'hb067, 16'ha80e, 16'ha180,
// 16'h9cdb, 16'h9a3a, 16'h99a6, 16'h9b2a,
// 16'h9eb0, 16'ha43c, 16'hab97, 16'hb4b1,
// 16'hbf4e, 16'hcb39, 16'hd83b, 16'he605,
// 16'hf45c, 16'h02ea, 16'h116c, 16'h1f93,
// 16'h2d17, 16'h39ae, 16'h451e, 16'h4f23,
// 16'h5792, 16'h5e37, 16'h62f7, 16'h65ae,
// 16'h6663, 16'h64f3, 16'h6189, 16'h5c19,
// 16'h54ce, 16'h4bd2, 16'h413e, 16'h3568,
// 16'h2871, 16'h1ab0, 16'h0c5c, 16'hfdd3,
// 16'hef48, 16'he123, 16'hd38f, 16'hc6ee,
// 16'hbb6b, 16'hb154, 16'ha8d1, 16'ha210,
// 16'h9d3e, 16'h9a63, 16'h999f, 16'h9aea,
// 16'h9e41, 16'ha395, 16'haac9, 16'hb3b4,
// 16'hbe2f, 16'hc9fb, 16'hd6e3, 16'he49c,
// 16'hf2eb, 16'h0172, 16'h0fff, 16'h1e2d,
// 16'h2bc6, 16'h3879, 16'h4407, 16'h4e37,
// 16'h56cb, 16'h5da5, 16'h6291, 16'h6584,
// 16'h6665, 16'h6532, 16'h61f7, 16'h5cba,
// 16'h559f, 16'h4cc7, 16'h4260, 16'h36a3,
// 16'h29c9, 16'h1c15, 16'h0dd2, 16'hff45,
// 16'hf0bc, 16'he286, 16'hd4e1, 16'hc826,
// 16'hbc81, 16'hb248, 16'ha992, 16'ha2ae,
// 16'h9d9d, 16'h9a99, 16'h9997, 16'h9ab3,
// 16'h9dd2, 16'ha2fa, 16'ha9fa, 16'hb2bd,
// 16'hbd13, 16'hc8be, 16'hd58e, 16'he338,
// 16'hf174, 16'h2002, 16'h0e88, 16'h1ccb,
// 16'h2a71, 16'h3742, 16'h42ee, 16'h4d42,
// 16'h5605, 16'h5d07, 16'h622e, 16'h654d,
// 16'h6669, 16'h6567, 16'h6261, 16'h5d56,
// 16'h5669, 16'h4dbd, 16'h437b, 16'h37de,
// 16'h2b1b, 16'h1d7e, 16'h0f40, 16'h20be,
// 16'hf22c, 16'he3ec, 16'hd637, 16'hc95e,
// 16'hbd9e, 16'hb33a, 16'haa61, 16'ha344,
// 16'h9e0d, 16'h9acb, 16'h999c, 16'h9a7d,
// 16'h9d6c, 16'ha25f, 16'ha931, 16'hb1cd,
// 16'hbbf6, 16'hc78a, 16'hd438, 16'he1d3,
// 16'hf003, 16'hfe8b, 16'h0d19, 16'h1b60,
// 16'h2920, 16'h3602, 16'h41d5, 16'h4c48,
// 16'h553a, 16'h5c69, 16'h61bf, 16'h6517,
// 16'h6661, 16'h659c, 16'h62c4, 16'h5dee,
// 16'h572f, 16'h4eaf, 16'h4491, 16'h3915,
// 16'h2c6e, 16'h1ee1, 16'h10b4, 16'h0231,
// 16'hf3a0, 16'he552, 16'hd78f, 16'hca99,
// 16'hbebf, 16'hb431, 16'hab30, 16'ha3e8,
// 16'h9e78, 16'h9b09, 16'h99a2, 16'h9a4d,
// 16'h9d0d, 16'ha1c7, 16'ha86f, 16'hb0dd,
// 16'hbae1, 16'hc653, 16'hd2e8, 16'he06f,
// 16'hee93, 16'hfd16, 16'h0ba4, 16'h19fb,
// 16'h27c5, 16'h34c6, 16'h40b4, 16'h4b4d,
// 16'h546a, 16'h5bc4, 16'h614f, 16'h64d6,
// 16'h665a, 16'h65c7, 16'h6324, 16'h5e80,
// 16'h57f2, 16'h4f98, 16'h45aa, 16'h3a45,
// 16'h2dc2, 16'h203f, 16'h1228, 16'h03a3,
// 16'hf515, 16'he6bd, 16'hd8e3, 16'hcbdd,
// 16'hbfdd, 16'hb530, 16'hac04, 16'ha48c,
// 16'h9eee, 16'h9b49, 16'h99ad, 16'h9a27,
// 16'h9cac, 16'ha13a, 16'ha7ae, 16'haff1,
// 16'hb9d2, 16'hc51d, 16'hd19c, 16'hdf0c,
// 16'hed22, 16'hfba1, 16'h0a33, 16'h188d,
// 16'h2670, 16'h3382, 16'h3f90, 16'h4a51,
// 16'h5390, 16'h5b21, 16'h60d4, 16'h6495,
// 16'h664a, 16'h65ee, 16'h637e, 16'h5f10,
// 16'h58ab, 16'h5086, 16'h46b5, 16'h3b7b,
// 16'h2f0a, 16'h21a6, 16'h1393, 16'h051c,
// 16'hf686, 16'he827, 16'hda3f, 16'hcd1e,
// 16'hc105, 16'hb62e, 16'hacdd, 16'ha535,
// 16'h9f69, 16'h9b8f, 16'h99bf, 16'h9a01,
// 16'h9c56, 16'ha0ac, 16'ha6f7, 16'haf08,
// 16'hb8c5, 16'hc3ec, 16'hd051, 16'hddaa,
// 16'hebb5, 16'hfa2c, 16'h08be, 16'h1723,
// 16'h2515, 16'h323c, 16'h3e6c, 16'h494d,
// 16'h52b7, 16'h5a73, 16'h6059, 16'h644a,
// 16'h663b, 16'h6609, 16'h63db, 16'h5f90,
// 16'h596b, 16'h5166, 16'h47c3, 16'h3ca9,
// 16'h3056, 16'h2304, 16'h1503, 16'h068e,
// 16'hf7fc, 16'he993, 16'hdb9c, 16'hce61,
// 16'hc22f, 16'hb731, 16'hadbb, 16'ha5e3,
// 16'h9fe8, 16'h9bd9, 16'h99d8, 16'h99e0,
// 16'h9c04, 16'ha027, 16'ha63e, 16'hae2a,
// 16'hb7b6, 16'hc2c2, 16'hcf06, 16'hdc4d,
// 16'hea46, 16'hf8b7, 16'h074a, 16'h15b7,
// 16'h23b7, 16'h30f7, 16'h3d40, 16'h4847,
// 16'h51d9, 16'h59c2, 16'h5fd6, 16'h6401,
// 16'h661a, 16'h662d, 16'h6424, 16'h601b,
// 16'h5a19, 16'h524a, 16'h48ca, 16'h3dd5,
// 16'h319c, 16'h2465, 16'h166e, 16'h0804,
// 16'hf971, 16'heafd, 16'hdcfc, 16'hcfab,
// 16'hc356, 16'hb83f, 16'hae96, 16'ha69b,
// 16'ha069, 16'h9c2b, 16'h99f3, 16'h99c7,
// 16'h9bb7, 16'h9fa4, 16'ha58f, 16'had49,
// 16'hb6b0, 16'hc19b, 16'hcdbc, 16'hdaf2,
// 16'he8d8, 16'hf743, 16'h05d6, 16'h1449,
// 16'h2257, 16'h2fb0, 16'h3c11, 16'h473f,
// 16'h50f4, 16'h590c, 16'h5f52, 16'h63ac,
// 16'h65fd, 16'h6642, 16'h6471, 16'h6097,
// 16'h5acb, 16'h5323, 16'h49d1, 16'h3efc,
// 16'h32e3, 16'h25bf, 16'h17db, 16'h0978,
// 16'hfae5, 16'hec6d, 16'hde5a, 16'hd0f6,
// 16'hc485, 16'hb94a, 16'haf7c, 16'ha753,
// 16'ha0f2, 16'h9c80, 16'h9a13, 16'h99b6,
// 16'h9b6b, 16'h9f2b, 16'ha4e0, 16'hac6f,
// 16'hb5b0, 16'hc070, 16'hcc7c, 16'hd993,
// 16'he76f, 16'hf5d0, 16'h045e, 16'h12dd,
// 16'h20f6, 16'h2e62, 16'h3ae5, 16'h462b,
// 16'h5013, 16'h584e, 16'h5ec9, 16'h6351,
// 16'h65dc, 16'h6652, 16'h64b7, 16'h6111,
// 16'h5b75, 16'h53fc, 16'h4ad1, 16'h4021,
// 16'h3425, 16'h271a, 16'h1946, 16'h0aea,
// 16'hfc5b, 16'hedde, 16'hdfb8, 16'hd247,
// 16'hc5b2, 16'hba5e, 16'hb063, 16'ha811,
// 16'ha17e, 16'h9cdc, 16'h9a39, 16'h99a8,
// 16'h9b27, 16'h9eb4, 16'ha438, 16'hab9a,
// 16'hb4b1, 16'hbf4b, 16'hcb3e, 16'hd835,
// 16'he60c, 16'hf456, 16'h02ef, 16'h1168,
// 16'h1f97, 16'h2d12, 16'h39b3, 16'h451b,
// 16'h4f24, 16'h5792, 16'h5e37, 16'h62f6,
// 16'h65b1, 16'h665e, 16'h64f8, 16'h6187,
// 16'h5c19, 16'h54cf, 16'h4bd0, 16'h413f,
// 16'h356b, 16'h286c, 16'h1ab3, 16'h0c5c,
// 16'hfdd0, 16'hef4d, 16'he11f, 16'hd390,
// 16'hc6ee, 16'hbb6b, 16'hb154, 16'ha8d0,
// 16'ha213, 16'h9d3a, 16'h9a67, 16'h999c,
// 16'h9ae9, 16'h9e45, 16'ha392, 16'haacb,
// 16'hb3b3, 16'hbe2e, 16'hc9fd, 16'hd6e0,
// 16'he4a1, 16'hf2e5, 16'h0178, 16'h0ffa,
// 16'h1e2f, 16'h2bc6, 16'h3878, 16'h440a,
// 16'h4e32, 16'h56d1, 16'h5d9e, 16'h6298,
// 16'h657e, 16'h6669, 16'h6531, 16'h61f6,
// 16'h5cbb, 16'h559d, 16'h4cc9, 16'h4261,
// 16'h36a1, 16'h29ca, 16'h1c14, 16'h0dd3,
// 16'hff44, 16'hf0bd, 16'he285, 16'hd4e2,
// 16'hc826, 16'hbc81, 16'hb245, 16'ha997,
// 16'ha2a9, 16'h9da0, 16'h9a98, 16'h9997,
// 16'h9ab4, 16'h9dd1, 16'ha2fb, 16'ha9f7,
// 16'hb2c3, 16'hbd0d, 16'hc8c1, 16'hd58f,
// 16'he335, 16'hf177, 16'hffff, 16'h0e8a,
// 16'h1ccb, 16'h2a71, 16'h3741, 16'h42ed,
// 16'h4d44, 16'h5604, 16'h5d0a, 16'h622a,
// 16'h6550, 16'h6665, 16'h656b, 16'h625f,
// 16'h5d56, 16'h566b, 16'h4db9, 16'h4380,
// 16'h37d9, 16'h2b1f, 16'h1d7a, 16'h0f44,
// 16'h20bb, 16'hf22f, 16'he3ea, 16'hd637,
// 16'hc95e, 16'hbd9f, 16'hb338, 16'haa64,
// 16'ha342, 16'h9e0e, 16'h9aca, 16'h999c,
// 16'h9a7d, 16'h9d6e, 16'ha25d, 16'ha932,
// 16'hb1cd, 16'hbbf4, 16'hc78d, 16'hd435,
// 16'he1d5, 16'hf002, 16'hfe8b, 16'h0d1a,
// 16'h1b5f, 16'h2920, 16'h3603, 16'h41d2,
// 16'h4c4d, 16'h5535, 16'h5c6d, 16'h61bd,
// 16'h6517, 16'h6662, 16'h659b, 16'h62c5,
// 16'h5ded, 16'h5730, 16'h4eae, 16'h4492,
// 16'h3916, 16'h2c6c, 16'h1ee3, 16'h10b2,
// 16'h0233, 16'hf39e, 16'he555, 16'hd78b,
// 16'hca9d, 16'hbebc, 16'hb433, 16'hab2f,
// 16'ha3e7, 16'h9e7a, 16'h9b08, 16'h99a3,
// 16'h9a4d, 16'h9d0c, 16'ha1c7, 16'ha871,
// 16'hb0da, 16'hbae5, 16'hc64f, 16'hd2ec,
// 16'he06b, 16'hee96, 16'hfd13, 16'h0ba8,
// 16'h19f7, 16'h27c8, 16'h34c5, 16'h40b2,
// 16'h4b51, 16'h5465, 16'h5bc9, 16'h614b,
// 16'h64da, 16'h6656, 16'h65cb, 16'h6320,
// 16'h5e84, 16'h57ee, 16'h4f9d, 16'h45a4,
// 16'h3a4c, 16'h2dba, 16'h2047, 16'h1222,
// 16'h03a7, 16'hf514, 16'he6bb, 16'hd8e6,
// 16'hcbdb, 16'hbfdf, 16'hb52f, 16'hac04,
// 16'ha48b, 16'h9ef0, 16'h9b48, 16'h99ae,
// 16'h9a26, 16'h9cad, 16'ha139, 16'ha7af,
// 16'haff1, 16'hb9d1, 16'hc51f, 16'hd19b,
// 16'hdf0b, 16'hed24, 16'hfba0, 16'h0a32,
// 16'h1890, 16'h266c, 16'h3385, 16'h3f90,
// 16'h4a4f, 16'h5393, 16'h5b1e, 16'h60d6,
// 16'h6494, 16'h664c, 16'h65eb, 16'h6382,
// 16'h5f0b, 16'h58b0, 16'h5083, 16'h46b5,
// 16'h3b7d, 16'h2f07, 16'h21a8, 16'h1393,
// 16'h0519, 16'hf68b, 16'he822, 16'hda43,
// 16'hcd1c, 16'hc105, 16'hb62f, 16'hacdb,
// 16'ha538, 16'h9f67, 16'h9b90, 16'h99bf,
// 16'h9a20, 16'h9c56, 16'ha0ae, 16'ha6f5,
// 16'haf0a, 16'hb8c2, 16'hc3ee, 16'hd051,
// 16'hdda9, 16'hebb8, 16'hfa27, 16'h08c2,
// 16'h1721, 16'h2515, 16'h323e, 16'h3e6a,
// 16'h494d, 16'h52b8, 16'h5a72, 16'h605a,
// 16'h644b, 16'h6637, 16'h660e, 16'h63d5,
// 16'h5f98, 16'h5963, 16'h516c, 16'h47bf,
// 16'h3cab, 16'h3055, 16'h2304, 16'h1504,
// 16'h068d, 16'hf7fd, 16'he993, 16'hdb9a,
// 16'hce65, 16'hc22b, 16'hb733, 16'hadbc,
// 16'ha5e1, 16'h9fe9, 16'h9bda, 16'h99d4,
// 16'h99e6, 16'h9bff, 16'ha029, 16'ha63f,
// 16'hae26, 16'hb7ba, 16'hc2c1, 16'hcf06,
// 16'hdc4c, 16'hea47, 16'hf8b6, 16'h074b,
// 16'h15b7, 16'h23b5, 16'h30fa, 16'h3d3e,
// 16'h4849, 16'h51d7, 16'h59c2, 16'h5fd9,
// 16'h63fc, 16'h661f, 16'h6629, 16'h6427,
// 16'h6018, 16'h5a1c, 16'h5247, 16'h48cc,
// 16'h3dd4, 16'h319d, 16'h2464, 16'h166e,
// 16'h0805, 16'hf970, 16'heaff, 16'hdcfa,
// 16'hcfab, 16'hc357, 16'hb83e, 16'hae98,
// 16'ha699, 16'ha069, 16'h9c2d, 16'h99ef,
// 16'h99cc, 16'h9bb2, 16'h9fa8, 16'ha58c,
// 16'had4a, 16'hb6b3, 16'hc193, 16'hcdc7,
// 16'hdae5, 16'he8e5, 16'hf73a, 16'h05db,
// 16'h1446, 16'h2259, 16'h2faf, 16'h3c12,
// 16'h473e, 16'h50f4, 16'h590d, 16'h5f51,
// 16'h63ac, 16'h65fe, 16'h6641, 16'h6471,
// 16'h6098, 16'h5aca, 16'h5323, 16'h49d2,
// 16'h3efa, 16'h32e5, 16'h25be, 16'h17db,
// 16'h0978, 16'hfae6, 16'hec6c, 16'hde5a,
// 16'hd0f6, 16'hc485, 16'hb94c, 16'haf7a,
// 16'ha753, 16'ha0f2, 16'h9c80, 16'h9a14,
// 16'h99b5, 16'h9b6b, 16'h9f2c, 16'ha4df,
// 16'hac70, 16'hb5ae, 16'hc072, 16'hcc7b,
// 16'hd994, 16'he76f, 16'hf5d0, 16'h045d,
// 16'h12df, 16'h20f3, 16'h2e65, 16'h3ae3,
// 16'h462d, 16'h5011, 16'h5850, 16'h5ec6,
// 16'h6355, 16'h65d8, 16'h6655, 16'h64b5,
// 16'h6113, 16'h5b73, 16'h53fd, 16'h4ad0,
// 16'h4022, 16'h3425, 16'h271a, 16'h1945,
// 16'h0aeb, 16'hfc5c, 16'heddb, 16'hdfbb,
// 16'hd244, 16'hc5b6, 16'hba5b, 16'hb064,
// 16'ha810, 16'ha180, 16'h9cdb, 16'h9a39,
// 16'h99a8, 16'h9b26, 16'h9eb7, 16'ha435,
// 16'hab9b, 16'hb4b0, 16'hbf4d, 16'hcb3c,
// 16'hd837, 16'he609, 16'hf458, 16'h02ed,
// 16'h116b, 16'h1f93, 16'h2d17, 16'h39ad,
// 16'h4520, 16'h4f20, 16'h5796, 16'h5e34,
// 16'h62f7, 16'h65b1, 16'h665d, 16'h64fa,
// 16'h6185, 16'h5c1a, 16'h54cf, 16'h4bcf,
// 16'h4141, 16'h3567, 16'h2872, 16'h1aad,
// 16'h0c60, 16'hfdce, 16'hef4e, 16'he11e,
// 16'hd391, 16'hc6ee, 16'hbb69, 16'hb158,
// 16'ha8cb, 16'ha216, 16'h9d3a, 16'h9a65,
// 16'h999e, 16'h9ae9, 16'h9e42, 16'ha396,
// 16'haac7, 16'hb3b6, 16'hbe2c, 16'hc9fe,
// 16'hd6e0, 16'he4a0, 16'hf2e7, 16'h0174,
// 16'h0fff, 16'h1e2b, 16'h2bc9, 16'h3876,
// 16'h440a, 16'h4e34, 16'h56ce, 16'h5da2,
// 16'h6293, 16'h6583, 16'h6665, 16'h6534,
// 16'h61f3, 16'h5cbf, 16'h559a, 16'h4ccb,
// 16'h425e, 16'h36a4, 16'h29c8, 16'h1c17,
// 16'h0dd0, 16'hff46, 16'hf0bc, 16'he284,
// 16'hd4e5, 16'hc822, 16'hbc86, 16'hb240,
// 16'ha99b, 16'ha2a5, 16'h9da6, 16'h9a90,
// 16'h99a0, 16'h9aab, 16'h9dd9, 16'ha2f5,
// 16'ha9fb, 16'hb2bf, 16'hbd11, 16'hc8bf,
// 16'hd58f, 16'he334, 16'hf179, 16'hfffe,
// 16'h0e8b, 16'h1cca, 16'h2a70, 16'h3743,
// 16'h42ed, 16'h4d43, 16'h5604, 16'h5d0b,
// 16'h6228, 16'h6552, 16'h6664, 16'h656c,
// 16'h625e, 16'h5d57, 16'h566a, 16'h4dbb,
// 16'h437e, 16'h37da, 16'h2b1f, 16'h1d7a,
// 16'h0f45, 16'h20b9, 16'hf230, 16'he3ea,
// 16'hd637, 16'hc95e, 16'hbd9e, 16'hb33a,
// 16'haa61, 16'ha346, 16'h9e09, 16'h9acf,
// 16'h9998, 16'h9a80, 16'h9d6c, 16'ha25d,
// 16'ha934, 16'hb1c9, 16'hbbfa, 16'hc787,
// 16'hd439, 16'he1d4, 16'hf020, 16'hfe8f,
// 16'h0d15, 16'h1b64, 16'h291c, 16'h3606,
// 16'h41d1, 16'h4c4c, 16'h5536, 16'h5c6d,
// 16'h61bb, 16'h651b, 16'h665e, 16'h659d,
// 16'h62c4, 16'h5dee, 16'h572f, 16'h4eaf,
// 16'h4490, 16'h3917, 16'h2c6d, 16'h1ee1,
// 16'h10b4, 16'h0230, 16'hf3a1, 16'he554,
// 16'hd78b, 16'hca9c, 16'hbebd, 16'hb432,
// 16'hab32, 16'ha3e3, 16'h9e7d, 16'h9b06,
// 16'h99a3, 16'h9a4f, 16'h9d09, 16'ha1ca,
// 16'ha86e, 16'hb0dc, 16'hbae4, 16'hc64f,
// 16'hd2eb, 16'he06e, 16'hee92, 16'hfd18,
// 16'h0ba2, 16'h19fb, 16'h27c7, 16'h34c4,
// 16'h40b5, 16'h4b4d, 16'h5468, 16'h5bc8,
// 16'h614a, 16'h64db, 16'h6657, 16'h65c7,
// 16'h6326, 16'h5e7e, 16'h57f4, 16'h4f97,
// 16'h45a8, 16'h3a49, 16'h2dbc, 16'h2047,
// 16'h1221, 16'h03a7, 16'hf513, 16'he6bc,
// 16'hd8e6, 16'hcbda, 16'hbfe0, 16'hb52d,
// 16'hac06, 16'ha48a, 16'h9ef0, 16'h9b48,
// 16'h99af, 16'h9a24, 16'h9caf, 16'ha137,
// 16'ha7b0, 16'haff3, 16'hb9ce, 16'hc522,
// 16'hd197, 16'hdf0f, 16'hed20, 16'hfba5,
// 16'h0a2d, 16'h1893, 16'h266c, 16'h3383,
// 16'h3f92, 16'h4a4e, 16'h5392, 16'h5b20,
// 16'h60d4, 16'h6496, 16'h6649, 16'h65ef,
// 16'h637d, 16'h5f10, 16'h58ac, 16'h5085,
// 16'h46b6, 16'h3b7a, 16'h2f0b, 16'h21a5,
// 16'h1395, 16'h0518, 16'hf68a, 16'he825,
// 16'hda40, 16'hcd1f, 16'hc101, 16'hb632,
// 16'hacda, 16'ha538, 16'h9f67, 16'h9b90,
// 16'h99bd, 16'h9a04, 16'h9c52, 16'ha0b1,
// 16'ha6f2, 16'haf0b, 16'hb8c4, 16'hc3eb,
// 16'hd054, 16'hdda6, 16'hebb9, 16'hfa28,
// 16'h08c0, 16'h1724, 16'h2511, 16'h3242,
// 16'h3e67, 16'h494f, 16'h52b7, 16'h5a71,
// 16'h605c, 16'h6449, 16'h6639, 16'h660c,
// 16'h63d8, 16'h5f93, 16'h596a, 16'h5164,
// 16'h47c6, 16'h3ca6, 16'h3058, 16'h2303,
// 16'h1505, 16'h068b, 16'hf820, 16'he98e,
// 16'hdb9f, 16'hce62, 16'hc22c, 16'hb735,
// 16'hadb7, 16'ha5e6, 16'h9fe6, 16'h9bdb,
// 16'h99d6, 16'h99e2, 16'h9c03, 16'ha026,
// 16'ha640, 16'hae27, 16'hb7b9, 16'hc2c0,
// 16'hcf09, 16'hdc47, 16'hea4c, 16'hf8b3,
// 16'h074c, 16'h15b7, 16'h23b5, 16'h30fa,
// 16'h3d3e, 16'h4848, 16'h51d8, 16'h59c2,
// 16'h5fd7, 16'h6420, 16'h661c, 16'h6629,
// 16'h642a, 16'h6013, 16'h5a21, 16'h5244,
// 16'h48cc, 16'h3dd7, 16'h3199, 16'h2467,
// 16'h166c, 16'h0805, 16'hf971, 16'heafd,
// 16'hdcfc, 16'hcfab, 16'hc356, 16'hb83f,
// 16'hae96, 16'ha69b, 16'ha06a, 16'h9c2a,
// 16'h99f2, 16'h99ca, 16'h9bb4, 16'h9fa7,
// 16'ha58c, 16'had4a, 16'hb6b1, 16'hc19a,
// 16'hcdbd, 16'hdaf0, 16'he8da, 16'hf743,
// 16'h05d5, 16'h144a, 16'h2256, 16'h2fb0,
// 16'h3c12, 16'h473d, 16'h50f7, 16'h5909,
// 16'h5f54, 16'h63a9, 16'h6601, 16'h663f,
// 16'h6473, 16'h6095, 16'h5acd, 16'h5322,
// 16'h49d1, 16'h3efd, 16'h32e0, 16'h25c4,
// 16'h17d6, 16'h097b, 16'hfae3, 16'hec6f,
// 16'hde59, 16'hd0f6, 16'hc486, 16'hb948,
// 16'haf7e, 16'ha751, 16'ha0f3, 16'h9c81,
// 16'h9a12, 16'h99b6, 16'h9b6b, 16'h9f2b,
// 16'ha4e0, 16'hac70, 16'hb5ae, 16'hc072,
// 16'hcc7b, 16'hd993, 16'he770, 16'hf5cf,
// 16'h045f, 16'h12dc, 16'h20f7, 16'h2e60,
// 16'h3ae8, 16'h4629, 16'h5014, 16'h584d,
// 16'h5eca, 16'h6350, 16'h65dd, 16'h6651,
// 16'h64b7, 16'h6112, 16'h5b73, 16'h53fe,
// 16'h4acf, 16'h4023, 16'h3423, 16'h271c,
// 16'h1944, 16'h0aec, 16'hfc5a, 16'heddd,
// 16'hdfba, 16'hd245, 16'hc5b4, 16'hba5d,
// 16'hb063, 16'ha810, 16'ha180, 16'h9cda,
// 16'h9a3b, 16'h99a6, 16'h9b28, 16'h9eb4,
// 16'ha438, 16'hab99, 16'hb4b1, 16'hbf4d,
// 16'hcb3b, 16'hd839, 16'he607, 16'hf45a,
// 16'h02ec, 16'h116b, 16'h1f93, 16'h2d17,
// 16'h39ae, 16'h451e, 16'h4f24, 16'h5791,
// 16'h5e36, 16'h62f8, 16'h65ae, 16'h6662,
// 16'h64f5, 16'h6188, 16'h5c17, 16'h54d3,
// 16'h4bcb, 16'h4144, 16'h3566, 16'h2871,
// 16'h1aaf, 16'h0c5f, 16'hfdce, 16'hef4e,
// 16'he11e, 16'hd392, 16'hc6ec, 16'hbb6d,
// 16'hb152, 16'ha8d1, 16'ha212, 16'h9d3c,
// 16'h9a64, 16'h999e, 16'h9aeb, 16'h9e3f,
// 16'ha399, 16'haac4, 16'hb3b9, 16'hbe2b,
// 16'hc9fe, 16'hd6e0, 16'he4a0, 16'hf2e7,
// 16'h0176, 16'h0ffc, 16'h1e2e, 16'h2bc5,
// 16'h387b, 16'h4406, 16'h4e36, 16'h56ce,
// 16'h5da0, 16'h6296, 16'h6581, 16'h6665,
// 16'h6535, 16'h61f2, 16'h5cbe, 16'h559c,
// 16'h4cca, 16'h425e, 16'h36a4, 16'h29c8,
// 16'h1c15, 16'h0dd3, 16'hff43, 16'hf0c0,
// 16'he281, 16'hd4e6, 16'hc820, 16'hbc87,
// 16'hb243, 16'ha997, 16'ha2a9, 16'h9da0,
// 16'h9a96, 16'h999b, 16'h9aaf, 16'h9dd7,
// 16'ha2f5, 16'ha9fc, 16'hb2be, 16'hbd11,
// 16'hc8c0, 16'hd58e, 16'he335, 16'hf179,
// 16'hfffc, 16'h0e8f, 16'h1cc4, 16'h2a77,
// 16'h373d, 16'h42f1, 16'h4d40, 16'h5607,
// 16'h5d07, 16'h622d, 16'h654d, 16'h6669,
// 16'h6568, 16'h6260, 16'h5d56, 16'h566b,
// 16'h4dba, 16'h437f, 16'h37d9, 16'h2b1f,
// 16'h1d7b, 16'h0f43, 16'h20bc, 16'hf22d,
// 16'he3ec, 16'hd635, 16'hc960, 16'hbd9e,
// 16'hb33a, 16'haa5f, 16'ha349, 16'h9e07,
// 16'h9ad0, 16'h9999, 16'h9a7d, 16'h9d6f,
// 16'ha25b, 16'ha935, 16'hb1c9, 16'hbbfa,
// 16'hc786, 16'hd43a, 16'he1d2, 16'hf004,
// 16'hfe8b, 16'h0d18, 16'h1b62, 16'h291e,
// 16'h3603, 16'h41d3, 16'h4c4b, 16'h5538,
// 16'h5c6c, 16'h61bb, 16'h6519, 16'h6660,
// 16'h659e, 16'h62c2, 16'h5def, 16'h572f,
// 16'h4eae, 16'h4492, 16'h3916, 16'h2c6c,
// 16'h1ee3, 16'h10b2, 16'h0232, 16'hf39f,
// 16'he555, 16'hd78b, 16'hca9c, 16'hbebd,
// 16'hb432, 16'hab30, 16'ha3e7, 16'h9e7a,
// 16'h9b07, 16'h99a4, 16'h9a4c, 16'h9d0d,
// 16'ha1c7, 16'ha86f, 16'hb0dd, 16'hbae1,
// 16'hc653, 16'hd2e8, 16'he06e, 16'hee95,
// 16'hfd13, 16'h0ba8, 16'h19f7, 16'h27c9,
// 16'h34c3, 16'h40b5, 16'h4b4e, 16'h5468,
// 16'h5bc7, 16'h614c, 16'h64d8, 16'h665a,
// 16'h65c5, 16'h6327, 16'h5e7e, 16'h57f2,
// 16'h4f9a, 16'h45a7, 16'h3a48, 16'h2dbf,
// 16'h2043, 16'h1224, 16'h03a7, 16'hf512,
// 16'he6bd, 16'hd8e5, 16'hcbdc, 16'hbfdd,
// 16'hb532, 16'hac20, 16'ha48f, 16'h9eed,
// 16'h9b49, 16'h99ae, 16'h9a26, 16'h9cac,
// 16'ha13b, 16'ha7ac, 16'haff4, 16'hb9cf,
// 16'hc51f, 16'hd19c, 16'hdf0a, 16'hed25,
// 16'hfb9f, 16'h0a33, 16'h188e, 16'h2670,
// 16'h3381, 16'h3f92, 16'h4a4e, 16'h5393,
// 16'h5b1f, 16'h60d5, 16'h6495, 16'h6649,
// 16'h65ef, 16'h637e, 16'h5f0e, 16'h58b0,
// 16'h507f, 16'h46bc, 16'h3b75, 16'h2f0e,
// 16'h21a5, 16'h1392, 16'h051c, 16'hf687,
// 16'he827, 16'hda3e, 16'hcd20, 16'hc101,
// 16'hb633, 16'hacd8, 16'ha53a, 16'h9f65,
// 16'h9b91, 16'h99bf, 16'h9a20, 16'h9c57,
// 16'ha0ac, 16'ha6f6, 16'haf0a, 16'hb8c2,
// 16'hc3ef, 16'hd04f, 16'hddab, 16'hebb5,
// 16'hfa2b, 16'h08be, 16'h1724, 16'h2513,
// 16'h323f, 16'h3e69, 16'h494f, 16'h52b5,
// 16'h5a74, 16'h605a, 16'h6449, 16'h663b,
// 16'h660a, 16'h63d8, 16'h5f94, 16'h5967,
// 16'h516a, 16'h47c0, 16'h3cac, 16'h3051,
// 16'h2309, 16'h14ff, 16'h0692, 16'hf7f9,
// 16'he994, 16'hdb9b, 16'hce63, 16'hc22d,
// 16'hb733, 16'hadb9, 16'ha5e5, 16'h9fe6,
// 16'h9bdc, 16'h99d5, 16'h99e2, 16'h9c03,
// 16'ha027, 16'ha63f, 16'hae29, 16'hb7b7,
// 16'hc2c1, 16'hcf07, 16'hdc4a, 16'hea4a,
// 16'hf8b5, 16'h074b, 16'h15b7, 16'h23b5,
// 16'h30f9, 16'h3d3f, 16'h4848, 16'h51d8,
// 16'h59c2, 16'h5fd7, 16'h63ff, 16'h661d,
// 16'h662a, 16'h6427, 16'h6017, 16'h5a1d,
// 16'h5246, 16'h48cd, 16'h3dd4, 16'h319d,
// 16'h2463, 16'h166f, 16'h0803, 16'hf972,
// 16'heafd, 16'hdcfc, 16'hcfa9, 16'hc35a,
// 16'hb83a, 16'hae9b, 16'ha697, 16'ha06c,
// 16'h9c2a, 16'h99f2, 16'h99c9, 16'h9bb4,
// 16'h9fa8, 16'ha58c, 16'had4a, 16'hb6b1,
// 16'hc197, 16'hcdc2, 16'hdaec, 16'he8dc,
// 16'hf742, 16'h05d5, 16'h144b, 16'h2255,
// 16'h2fb1, 16'h3c10, 16'h473f, 16'h50f6,
// 16'h590a, 16'h5f53, 16'h63aa, 16'h65ff,
// 16'h6642, 16'h646f, 16'h609a, 16'h5ac7,
// 16'h5328, 16'h49cc, 16'h3f20, 16'h32df,
// 16'h25c3, 16'h17d7, 16'h097b, 16'hfae3,
// 16'hec70, 16'hde56, 16'hd0fa, 16'hc481,
// 16'hb94d, 16'haf7c, 16'ha751, 16'ha0f4,
// 16'h9c7f, 16'h9a13, 16'h99b6, 16'h9b6c,
// 16'h9f2a, 16'ha4e1, 16'hac6e, 16'hb5b0,
// 16'hc071, 16'hcc7c, 16'hd992, 16'he772,
// 16'hf5cb, 16'h0464, 16'h12d8, 16'h20f8,
// 16'h2e63, 16'h3ae2, 16'h462f, 16'h500f,
// 16'h5851, 16'h5ec6, 16'h6355, 16'h65d7,
// 16'h6656, 16'h64b5, 16'h6111, 16'h5b76,
// 16'h53fa, 16'h4ad2, 16'h4023, 16'h3422,
// 16'h271d, 16'h1942, 16'h0aee, 16'hfc59,
// 16'heddd, 16'hdfbb, 16'hd243, 16'hc5b7,
// 16'hba59, 16'hb066, 16'ha80f, 16'ha17f,
// 16'h9cde, 16'h9a35, 16'h99ac, 16'h9b24,
// 16'h9eb6, 16'ha438, 16'hab99, 16'hb4b1,
// 16'hbf4c, 16'hcb3d, 16'hd837, 16'he608,
// 16'hf45a, 16'h02eb, 16'h116c, 16'h1f93,
// 16'h2d16, 16'h39af, 16'h451e, 16'h4f23,
// 16'h5792, 16'h5e37, 16'h62f6, 16'h65b0,
// 16'h6661, 16'h64f5, 16'h6188, 16'h5c19,
// 16'h54cf, 16'h4bce, 16'h4144, 16'h3563,
// 16'h2875, 16'h1aac, 16'h0c60, 16'hfdce,
// 16'hef4f, 16'he11c, 16'hd394, 16'hc6ea,
// 16'hbb6f, 16'hb152, 16'ha8d0, 16'ha213,
// 16'h9d39, 16'h9a69, 16'h999a, 16'h9aec,
// 16'h9e41, 16'ha395, 16'haaca, 16'hb3b2,
// 16'hbe30, 16'hc9fa, 16'hd6e5, 16'he49c,
// 16'hf2e9, 16'h0174, 16'h0ffd, 16'h1e2e,
// 16'h2bc6, 16'h3879, 16'h4407, 16'h4e36,
// 16'h56cd, 16'h5da2, 16'h6294, 16'h6581,
// 16'h6667, 16'h6533, 16'h61f4, 16'h5cbc,
// 16'h559e, 16'h4cc7, 16'h4262, 16'h36a1,
// 16'h29c9, 16'h1c16, 16'h0dd0, 16'hff48,
// 16'hf0ba, 16'he285, 16'hd4e4, 16'hc822,
// 16'hbc86, 16'hb243, 16'ha996, 16'ha2ab,
// 16'h9d9f, 16'h9a98, 16'h9997, 16'h9ab4,
// 16'h9dd3, 16'ha2f7, 16'ha9fc, 16'hb2bd,
// 16'hbd12, 16'hc8c0, 16'hd58d, 16'he336,
// 16'hf177, 16'h2020, 16'h0e89, 16'h1ccb,
// 16'h2a71, 16'h3741, 16'h42ef, 16'h4d41,
// 16'h5606, 16'h5d08, 16'h622c, 16'h654f,
// 16'h6667, 16'h6568, 16'h6262, 16'h5d53,
// 16'h566e, 16'h4db9, 16'h437d, 16'h37dc,
// 16'h2b1d, 16'h1d7c, 16'h0f43, 16'h20ba,
// 16'hf230, 16'he3e8, 16'hd63b, 16'hc959,
// 16'hbda4, 16'hb334, 16'haa66, 16'ha341,
// 16'h9e0f, 16'h9ac8, 16'h99a0, 16'h9a79,
// 16'h9d70, 16'ha25c, 16'ha933, 16'hb1cb,
// 16'hbbf8, 16'hc787, 16'hd43b, 16'he1d2,
// 16'hf002, 16'hfe8c, 16'h0d18, 16'h1b62,
// 16'h291e, 16'h3604, 16'h41d2, 16'h4c4b,
// 16'h5538, 16'h5c6a, 16'h61c0, 16'h6515,
// 16'h6663, 16'h659b, 16'h62c3, 16'h5def,
// 16'h5731, 16'h4eaa, 16'h4497, 16'h3911,
// 16'h2c6f, 16'h1ee2, 16'h10b3, 16'h0230,
// 16'hf3a2, 16'he551, 16'hd78e, 16'hca9c,
// 16'hbebb, 16'hb435, 16'hab2d, 16'ha3e9,
// 16'h9e78, 16'h9b0a, 16'h99a0, 16'h9a51,
// 16'h9d08, 16'ha1cb, 16'ha86e, 16'hb0da,
// 16'hbae6, 16'hc64e, 16'hd2ec, 16'he06c,
// 16'hee95, 16'hfd14, 16'h0ba6, 16'h19f8,
// 16'h27c8, 16'h34c5, 16'h40b3, 16'h4b4f,
// 16'h5467, 16'h5bc8, 16'h614a, 16'h64dc,
// 16'h6655, 16'h65c9, 16'h6324, 16'h5e7f,
// 16'h57f4, 16'h4f97, 16'h45a8, 16'h3a49,
// 16'h2dbd, 16'h2045, 16'h1222, 16'h03a7,
// 16'hf515, 16'he6ba, 16'hd8e7, 16'hcbda,
// 16'hbfdd, 16'hb533, 16'hac20, 16'ha48f,
// 16'h9eed, 16'h9b48, 16'h99b0, 16'h9a23,
// 16'h9caf, 16'ha137, 16'ha7b2, 16'hafed,
// 16'hb9d6, 16'hc51a, 16'hd19d, 16'hdf0b,
// 16'hed23, 16'hfba2, 16'h0a31, 16'h188f,
// 16'h266d, 16'h3385, 16'h3f8f, 16'h4a51,
// 16'h5391, 16'h5b1e, 16'h60d7, 16'h6493,
// 16'h664c, 16'h65ec, 16'h6381, 16'h5f0b,
// 16'h58b0, 16'h5083, 16'h46b6, 16'h3b7b,
// 16'h2f09, 16'h21a8, 16'h1392, 16'h051b,
// 16'hf687, 16'he826, 16'hda41, 16'hcd1d,
// 16'hc103, 16'hb631, 16'hacda, 16'ha539,
// 16'h9f66, 16'h9b8f, 16'h99c0, 16'h9a20,
// 16'h9c57, 16'ha0ad, 16'ha6f5, 16'haf0a,
// 16'hb8c3, 16'hc3ed, 16'hd052, 16'hdda8,
// 16'hebb8, 16'hfa28, 16'h08c1, 16'h1721,
// 16'h2515, 16'h323e, 16'h3e6a, 16'h494e,
// 16'h52b6, 16'h5a74, 16'h6057, 16'h644e,
// 16'h6636, 16'h660e, 16'h63d6, 16'h5f94,
// 16'h5968, 16'h5168, 16'h47c2, 16'h3caa,
// 16'h3053, 16'h2308, 16'h1520, 16'h068f,
// 16'hf7fd, 16'he992, 16'hdb9b, 16'hce65,
// 16'hc229, 16'hb737, 16'hadb7, 16'ha5e5,
// 16'h9fe8, 16'h9bd8, 16'h99d8, 16'h99e1,
// 16'h9c03, 16'ha027, 16'ha640, 16'hae26,
// 16'hb7b9, 16'hc2c2, 16'hcf05, 16'hdc4d,
// 16'hea46, 16'hf8b8, 16'h0748, 16'h15bb,
// 16'h23b1, 16'h30fc, 16'h3d3e, 16'h4847,
// 16'h51da, 16'h59bf, 16'h5fdb, 16'h63fa,
// 16'h6622, 16'h6626, 16'h6428, 16'h6019,
// 16'h5a1a, 16'h5248, 16'h48cd, 16'h3dd2,
// 16'h319f, 16'h2463, 16'h166d, 16'h0806,
// 16'hf970, 16'heafe, 16'hdcfb, 16'hcfaa,
// 16'hc358, 16'hb83d, 16'hae99, 16'ha697,
// 16'ha06d, 16'h9c27, 16'h99f6, 16'h99c6,
// 16'h9bb6, 16'h9fa7, 16'ha58b, 16'had4c,
// 16'hb6b0, 16'hc198, 16'hcdc0, 16'hdaee,
// 16'he8db, 16'hf743, 16'h05d4, 16'h144b,
// 16'h2257, 16'h2fad, 16'h3c16, 16'h4739,
// 16'h50fa, 16'h5908, 16'h5f54, 16'h63aa,
// 16'h65ff, 16'h6641, 16'h6471, 16'h6098,
// 16'h5ac9, 16'h5325, 16'h49cf, 16'h3efe,
// 16'h32e1, 16'h25c0, 16'h17db, 16'h0976,
// 16'hfae8, 16'hec6b, 16'hde5b, 16'hd0f6,
// 16'hc484, 16'hb94b, 16'haf7c, 16'ha753,
// 16'ha0f1, 16'h9c82, 16'h9a11, 16'h99b7,
// 16'h9b6b, 16'h9f2a, 16'ha4e2, 16'hac6d,
// 16'hb5b1, 16'hc070, 16'hcc7c, 16'hd992,
// 16'he772, 16'hf5cc, 16'h0463, 16'h12d9,
// 16'h20f6, 16'h2e65, 16'h3ae1, 16'h4630,
// 16'h500f, 16'h5850, 16'h5ec7, 16'h6353,
// 16'h65db, 16'h6652, 16'h64b7, 16'h6112,
// 16'h5b73, 16'h53fe, 16'h4ace, 16'h4024,
// 16'h3424, 16'h271a, 16'h1946, 16'h0aea,
// 16'hfc5c, 16'heddb, 16'hdfbc, 16'hd242,
// 16'hc5b8, 16'hba59, 16'hb067, 16'ha80c,
// 16'ha183, 16'h9cd9, 16'h9a3a, 16'h99a8,
// 16'h9b26, 16'h9eb6, 16'ha438, 16'hab98,
// 16'hb4b1, 16'hbf4e, 16'hcb39, 16'hd83c,
// 16'he604, 16'hf45d, 16'h02e9, 16'h116d,
// 16'h1f92, 16'h2d17, 16'h39af, 16'h451d,
// 16'h4f24, 16'h5792, 16'h5e35, 16'h62f9,
// 16'h65ae, 16'h6660, 16'h64f8, 16'h6185,
// 16'h5c1b, 16'h54ce, 16'h4bcf, 16'h4143,
// 16'h3565, 16'h2873, 16'h1aac, 16'h0c61,
// 16'hfdcf, 16'hef4d, 16'he11d, 16'hd394,
// 16'hc6ea, 16'hbb6f, 16'hb151, 16'ha8d2,
// 16'ha211, 16'h9d3c, 16'h9a65, 16'h999d,
// 16'h9aeb, 16'h9e41, 16'ha396, 16'haac7,
// 16'hb3b6, 16'hbe2d, 16'hc9fc, 16'hd6e4,
// 16'he49b, 16'hf2ea, 16'h0174, 16'h0ffd,
// 16'h1e2e, 16'h2bc6, 16'h3877, 16'h440b,
// 16'h4e32, 16'h56d0, 16'h5da0, 16'h6294,
// 16'h6584, 16'h6663, 16'h6535, 16'h61f4,
// 16'h5cbb, 16'h559f, 16'h4cc7, 16'h4261,
// 16'h36a2, 16'h29c9, 16'h1c16, 16'h0dd0,
// 16'hff47, 16'hf0bc, 16'he284, 16'hd4e4,
// 16'hc822, 16'hbc85, 16'hb244, 16'ha997,
// 16'ha2a8, 16'h9da2, 16'h9a95, 16'h999b,
// 16'h9aaf, 16'h9dd6, 16'ha2f7, 16'ha9fb,
// 16'hb2be, 16'hbd11, 16'hc8c0, 16'hd58d,
// 16'he338, 16'hf174, 16'h2002, 16'h0e88,
// 16'h1ccb, 16'h2a71, 16'h3743, 16'h42ec,
// 16'h4d43, 16'h5605, 16'h5d09, 16'h622b,
// 16'h6550, 16'h6665, 16'h656b, 16'h625f,
// 16'h5d56, 16'h566a, 16'h4dbd, 16'h437a,
// 16'h37de, 16'h2b1c, 16'h1d7c, 16'h0f44,
// 16'h20b9, 16'hf230, 16'he3ea, 16'hd637,
// 16'hc95e, 16'hbda0, 16'hb337, 16'haa63,
// 16'ha343, 16'h9e0d, 16'h9acc, 16'h999a,
// 16'h9a7f, 16'h9d6a, 16'ha261, 16'ha930,
// 16'hb1cd, 16'hbbf6, 16'hc789, 16'hd438,
// 16'he1d5, 16'hf001, 16'hfe8d, 16'h0d16,
// 16'h1b64, 16'h291c, 16'h3605, 16'h41d2,
// 16'h4c4b, 16'h5538, 16'h5c6b, 16'h61be,
// 16'h6515, 16'h6664, 16'h659a, 16'h62c4,
// 16'h5df0, 16'h572d, 16'h4eaf, 16'h4492,
// 16'h3914, 16'h2c6f, 16'h1ee0, 16'h10b5,
// 16'h022f, 16'hf3a2, 16'he552, 16'hd78d,
// 16'hca9b, 16'hbebe, 16'hb431, 16'hab32,
// 16'ha3e4, 16'h9e7c, 16'h9b07, 16'h99a3,
// 16'h9a4e, 16'h9d0a, 16'ha1ca, 16'ha86d,
// 16'hb0de, 16'hbae1, 16'hc652, 16'hd2ea,
// 16'he06d, 16'hee94, 16'hfd14, 16'h0ba7,
// 16'h19f8, 16'h27c8, 16'h34c5, 16'h40b2,
// 16'h4b50, 16'h5467, 16'h5bc7, 16'h614c,
// 16'h64d9, 16'h6657, 16'h65c9, 16'h6323,
// 16'h5e81, 16'h57f0, 16'h4f9c, 16'h45a5,
// 16'h3a4a, 16'h2dbc, 16'h2046, 16'h1222,
// 16'h03a9, 16'hf510, 16'he6bf, 16'hd8e2,
// 16'hcbdf, 16'hbfdc, 16'hb530, 16'hac03,
// 16'ha48c, 16'h9eef, 16'h9b49, 16'h99ae,
// 16'h9a23, 16'h9cb1, 16'ha134, 16'ha7b5,
// 16'hafeb, 16'hb9d7, 16'hc518, 16'hd1a2,
// 16'hdf06, 16'hed26, 16'hfba0, 16'h0a31,
// 16'h1891, 16'h266d, 16'h3383, 16'h3f91,
// 16'h4a4f, 16'h5392, 16'h5b1f, 16'h60d5,
// 16'h6496, 16'h6649, 16'h65ee, 16'h637e,
// 16'h5f10, 16'h58ab, 16'h5087, 16'h46b2,
// 16'h3b7f, 16'h2f07, 16'h21a8, 16'h1392,
// 16'h051b, 16'hf688, 16'he826, 16'hda3f,
// 16'hcd1f, 16'hc102, 16'hb632, 16'hacd9,
// 16'ha53a, 16'h9f63, 16'h9b94, 16'h99bb,
// 16'h9a04, 16'h9c55, 16'ha0ab, 16'ha6f9,
// 16'haf06, 16'hb8c6, 16'hc3ec, 16'hd051,
// 16'hddaa, 16'hebb5, 16'hfa2c, 16'h08bd,
// 16'h1725, 16'h2512, 16'h3240, 16'h3e69,
// 16'h494e, 16'h52b6, 16'h5a74, 16'h6058,
// 16'h644d, 16'h6636, 16'h660e, 16'h63d6,
// 16'h5f94, 16'h596a, 16'h5165, 16'h47c4,
// 16'h3ca8, 16'h3055, 16'h2307, 16'h1501,
// 16'h068e, 16'hf7fd, 16'he992, 16'hdb9b,
// 16'hce66, 16'hc228, 16'hb738, 16'hadb5,
// 16'ha5e8, 16'h9fe5, 16'h9bdb, 16'h99d5,
// 16'h99e4, 16'h9c20, 16'ha02b, 16'ha63a,
// 16'hae2c, 16'hb7b6, 16'hc2c1, 16'hcf08,
// 16'hdc4a, 16'hea48, 16'hf8b8, 16'h0747,
// 16'h15ba, 16'h23b4, 16'h30f9, 16'h3d41,
// 16'h4845, 16'h51db, 16'h59bf, 16'h5fd9,
// 16'h63ff, 16'h661b, 16'h662e, 16'h6422,
// 16'h601c, 16'h5a19, 16'h5249, 16'h48ca,
// 16'h3dd6, 16'h319b, 16'h2467, 16'h166a,
// 16'h0808, 16'hf96d, 16'heb02, 16'hdcf8,
// 16'hcfac, 16'hc357, 16'hb83e, 16'hae97,
// 16'ha69b, 16'ha067, 16'h9c2f, 16'h99ed,
// 16'h99ce, 16'h9bb0, 16'h9faa, 16'ha58c,
// 16'had48, 16'hb6b4, 16'hc194, 16'hcdc4,
// 16'hdaeb, 16'he8de, 16'hf73f, 16'h05d7,
// 16'h1449, 16'h2257, 16'h2fb0, 16'h3c12,
// 16'h473d, 16'h50f6, 16'h590a, 16'h5f54,
// 16'h63aa, 16'h65ff, 16'h6641, 16'h6470,
// 16'h6099, 16'h5ac9, 16'h5325, 16'h49d0,
// 16'h3efc, 16'h32e2, 16'h25c1, 16'h17d8,
// 16'h097c, 16'hfae1, 16'hec70, 16'hde58,
// 16'hd0f7, 16'hc484, 16'hb94c, 16'haf7a,
// 16'ha754, 16'ha0f2, 16'h9c7f, 16'h9a15,
// 16'h99b3, 16'h9b6e, 16'h9f29, 16'ha4e1,
// 16'hac6f, 16'hb5af, 16'hc070, 16'hcc7e,
// 16'hd98f, 16'he775, 16'hf5ca, 16'h0463,
// 16'h12d9, 16'h20f8, 16'h2e61, 16'h3ae6,
// 16'h462b, 16'h5012, 16'h584f, 16'h5ec8,
// 16'h6352, 16'h65db, 16'h6652, 16'h64b8,
// 16'h6110, 16'h5b75, 16'h53fc, 16'h4ad0,
// 16'h4022, 16'h3426, 16'h2718, 16'h1947,
// 16'h0aeb, 16'hfc58, 16'hede1, 16'hdfb7,
// 16'hd245, 16'hc5b7, 16'hba58, 16'hb068,
// 16'ha80e, 16'ha17f, 16'h9cdc, 16'h9a3a,
// 16'h99a6, 16'h9b29, 16'h9eb3, 16'ha438,
// 16'hab9b, 16'hb4af, 16'hbf4e, 16'hcb3b,
// 16'hd838, 16'he608, 16'hf45a, 16'h02eb,
// 16'h116d, 16'h1f91, 16'h2d18, 16'h39ad,
// 16'h451e, 16'h4f25, 16'h5790, 16'h5e39,
// 16'h62f3, 16'h65b3, 16'h665e, 16'h64f8,
// 16'h6186, 16'h5c19, 16'h54d0, 16'h4bcf,
// 16'h4141, 16'h3567, 16'h2871, 16'h1aae,
// 16'h0c5f, 16'hfdd0, 16'hef4c, 16'he11f,
// 16'hd392, 16'hc6eb, 16'hbb6e, 16'hb153,
// 16'ha8cf, 16'ha214, 16'h9d3a, 16'h9a66,
// 16'h999d, 16'h9aea, 16'h9e42, 16'ha396,
// 16'haac6, 16'hb3b7, 16'hbe2c, 16'hc9fe,
// 16'hd6e1, 16'he49e, 16'hf2e8, 16'h0176,
// 16'h0ffa, 16'h1e31, 16'h2bc3, 16'h387c,
// 16'h4405, 16'h4e37, 16'h56cc, 16'h5da4,
// 16'h6292, 16'h6584, 16'h6663, 16'h6536,
// 16'h61f3, 16'h5cbc, 16'h559e, 16'h4cc8,
// 16'h4260, 16'h36a3, 16'h29c7, 16'h1c17,
// 16'h0dd1, 16'hff45, 16'hf0bd, 16'he285,
// 16'hd4e1, 16'hc826, 16'hbc82, 16'hb245,
// 16'ha997, 16'ha2a9, 16'h9d9f, 16'h9a9a,
// 16'h9995, 16'h9ab5, 16'h9dd2, 16'ha2f8,
// 16'ha9fb, 16'hb2bf, 16'hbd0f, 16'hc8c3,
// 16'hd58a, 16'he339, 16'hf176, 16'hfffe,
// 16'h0e8c, 16'h1cc9, 16'h2a72, 16'h3741,
// 16'h42ee, 16'h4d42, 16'h5605, 16'h5d09,
// 16'h622c, 16'h654d, 16'h6669, 16'h6568,
// 16'h625f, 16'h5d5a, 16'h5664, 16'h4dc1,
// 16'h4379, 16'h37de, 16'h2b1d, 16'h1d7a,
// 16'h0f45, 16'h20b9, 16'hf231, 16'he3e8,
// 16'hd639, 16'hc95d, 16'hbd9f, 16'hb339,
// 16'haa61, 16'ha345, 16'h9e0d, 16'h9aca,
// 16'h999c, 16'h9a7e, 16'h9d6b, 16'ha260,
// 16'ha930, 16'hb1cd, 16'hbbf7, 16'hc789,
// 16'hd438, 16'he1d2, 16'hf005, 16'hfe89,
// 16'h0d1b, 16'h1b5f, 16'h2920, 16'h3602,
// 16'h41d4, 16'h4c4a, 16'h5539, 16'h5c69,
// 16'h61c0, 16'h6514, 16'h6665, 16'h6599,
// 16'h62c5, 16'h5dee, 16'h5730, 16'h4eac,
// 16'h4495, 16'h3912, 16'h2c6f, 16'h1ee2,
// 16'h10b2, 16'h0232, 16'hf3a0, 16'he552,
// 16'hd78f, 16'hca99, 16'hbebe, 16'hb432,
// 16'hab30, 16'ha3e7, 16'h9e79, 16'h9b09,
// 16'h99a1, 16'h9a4f, 16'h9d0b, 16'ha1c7,
// 16'ha871, 16'hb0da, 16'hbae4, 16'hc650,
// 16'hd2eb, 16'he06c, 16'hee96, 16'hfd12,
// 16'h0ba9, 16'h19f7, 16'h27c7, 16'h34c6,
// 16'h40b2, 16'h4b50, 16'h5467, 16'h5bc6,
// 16'h614e, 16'h64d7, 16'h6659, 16'h65c7,
// 16'h6324, 16'h5e81, 16'h57f1, 16'h4f9a,
// 16'h45a7, 16'h3a48, 16'h2dbe, 16'h2044,
// 16'h1224, 16'h03a7, 16'hf512, 16'he6bd,
// 16'hd8e4, 16'hcbdc, 16'hbfdf, 16'hb52f,
// 16'hac04, 16'ha48b, 16'h9eef, 16'h9b48,
// 16'h99b1, 16'h9a21, 16'h9cb1, 16'ha135,
// 16'ha7b3, 16'hafee, 16'hb9d4, 16'hc51a,
// 16'hd19f, 16'hdf09, 16'hed25, 16'hfba1,
// 16'h0a2f, 16'h1892, 16'h266d, 16'h3383,
// 16'h3f91, 16'h4a4f, 16'h5392, 16'h5b20,
// 16'h60d4, 16'h6495, 16'h664a, 16'h65ed,
// 16'h6381, 16'h5f0c, 16'h58af, 16'h5083,
// 16'h46b5, 16'h3b7c, 16'h2f0a, 16'h21a6,
// 16'h1394, 16'h0519, 16'hf688, 16'he827,
// 16'hda3f, 16'hcd1f, 16'hc103, 16'hb62f,
// 16'hacdd, 16'ha535, 16'h9f6a, 16'h9b8d,
// 16'h99c0, 16'h9a01, 16'h9c55, 16'ha0ae,
// 16'ha6f4, 16'haf0b, 16'hb8c1, 16'hc3f1,
// 16'hd04d, 16'hddac, 16'hebb4, 16'hfa2c,
// 16'h08be, 16'h1725, 16'h2511, 16'h3241,
// 16'h3e68, 16'h494f, 16'h52b5, 16'h5a75,
// 16'h6057, 16'h644f, 16'h6633, 16'h6611,
// 16'h63d3, 16'h5f97, 16'h5967, 16'h5167,
// 16'h47c3, 16'h3ca9, 16'h3054, 16'h2307,
// 16'h1520, 16'h0691, 16'hf7fb, 16'he991,
// 16'hdb9e, 16'hce60, 16'hc230, 16'hb731,
// 16'hadbb, 16'ha5e2, 16'h9fea, 16'h9bd7,
// 16'h99d9, 16'h99e1, 16'h9c02, 16'ha029,
// 16'ha63c, 16'hae2a, 16'hb7b8, 16'hc2c1,
// 16'hcf07, 16'hdc4a, 16'hea48, 16'hf8b7,
// 16'h0749, 16'h15ba, 16'h23b2, 16'h30fc,
// 16'h3d3d, 16'h4848, 16'h51d9, 16'h59c0,
// 16'h5fd9, 16'h63ff, 16'h661b, 16'h662d,
// 16'h6422, 16'h601d, 16'h5a18, 16'h524a,
// 16'h48ca, 16'h3dd5, 16'h319c, 16'h2465,
// 16'h166e, 16'h0804, 16'hf971, 16'heafd,
// 16'hdcfc, 16'hcfab, 16'hc357, 16'hb83e,
// 16'hae95, 16'ha69e, 16'ha066, 16'h9c2e,
// 16'h99ef, 16'h99cb, 16'h9bb4, 16'h9fa6,
// 16'ha58e, 16'had48, 16'hb6b4, 16'hc195,
// 16'hcdc2, 16'hdaec, 16'he8dd, 16'hf741,
// 16'h05d6, 16'h1449, 16'h2257, 16'h2fb0,
// 16'h3c11, 16'h473f, 16'h50f3, 16'h590e,
// 16'h5f50, 16'h63ac, 16'h65ff, 16'h6640,
// 16'h6472, 16'h6096, 16'h5acd, 16'h5320,
// 16'h49d5, 16'h3ef9, 16'h32e3, 16'h25c2,
// 16'h17d6, 16'h097d, 16'hfae2, 16'hec6e,
// 16'hde5b, 16'hd0f4, 16'hc487, 16'hb949,
// 16'haf7d, 16'ha752, 16'ha0f2, 16'h9c81,
// 16'h9a12, 16'h99b7, 16'h9b6a, 16'h9f2c,
// 16'ha4de, 16'hac73, 16'hb5aa, 16'hc076,
// 16'hcc78, 16'hd995, 16'he76f, 16'hf5ce,
// 16'h0462, 16'h12d9, 16'h20f8, 16'h2e62,
// 16'h3ae3, 16'h462f, 16'h500f, 16'h5850,
// 16'h5ec8, 16'h6352, 16'h65db, 16'h6652,
// 16'h64b7, 16'h6112, 16'h5b72, 16'h5420,
// 16'h4acc, 16'h4027, 16'h341f, 16'h271f,
// 16'h1941, 16'h0aef, 16'hfc58, 16'hedde,
// 16'hdfba, 16'hd244, 16'hc5b6, 16'hba59,
// 16'hb068, 16'ha80c, 16'ha182, 16'h9cdb,
// 16'h9a39, 16'h99a7, 16'h9b28, 16'h9eb3,
// 16'ha439, 16'hab9a, 16'hb4af, 16'hbf4f,
// 16'hcb38, 16'hd83c, 16'he605, 16'hf45b,
// 16'h02eb, 16'h116c, 16'h1f93, 16'h2d16,
// 16'h39b0, 16'h451b, 16'h4f26, 16'h5791,
// 16'h5e36, 16'h62f8, 16'h65af, 16'h665f,
// 16'h64f9, 16'h6183, 16'h5c1e, 16'h54cc,
// 16'h4bd1, 16'h4140, 16'h3568, 16'h2870,
// 16'h1aaf, 16'h0c60, 16'hfdcd, 16'hef50,
// 16'he11c, 16'hd392, 16'hc6ed, 16'hbb6c,
// 16'hb153, 16'ha8d2, 16'ha20f, 16'h9d3f,
// 16'h9a62, 16'h99a0, 16'h9ae9, 16'h9e41,
// 16'ha397, 16'haac6, 16'hb3b7, 16'hbe2d,
// 16'hc9fb, 16'hd6e4, 16'he49d, 16'hf2e7,
// 16'h0177, 16'h0ffb, 16'h1e2e, 16'h2bc8,
// 16'h3876, 16'h4409, 16'h4e35, 16'h56cd,
// 16'h5da4, 16'h6292, 16'h6582, 16'h6666,
// 16'h6533, 16'h61f6, 16'h5cba, 16'h559f,
// 16'h4cc7, 16'h4260, 16'h36a4, 16'h29c7,
// 16'h1c18, 16'h0dcf, 16'hff47, 16'hf0bb,
// 16'he286, 16'hd4e2, 16'hc824, 16'hbc84,
// 16'hb245, 16'ha994, 16'ha2ac, 16'h9d9d,
// 16'h9a9b, 16'h9995, 16'h9ab5, 16'h9dd0,
// 16'ha2fc, 16'ha9f7, 16'hb2c1, 16'hbd0f,
// 16'hc8c1, 16'hd58d, 16'he337, 16'hf176,
// 16'hffff, 16'h0e8b, 16'h1cc9, 16'h2a73,
// 16'h3740, 16'h42ef, 16'h4d42, 16'h5605,
// 16'h5d09, 16'h622a, 16'h6551, 16'h6666,
// 16'h6569, 16'h6260, 16'h5d56, 16'h5669,
// 16'h4dbe, 16'h4379, 16'h37df, 16'h2b1b,
// 16'h1d7d, 16'h0f42, 16'h20bc, 16'hf22d,
// 16'he3ed, 16'hd634, 16'hc961, 16'hbd9c,
// 16'hb33b, 16'haa61, 16'ha344, 16'h9e0d,
// 16'h9acb, 16'h999c, 16'h9a7d, 16'h9d6c,
// 16'ha25f, 16'ha932, 16'hb1cb, 16'hbbf9,
// 16'hc785, 16'hd43d, 16'he1cf, 16'hf006,
// 16'hfe89, 16'h0d19, 16'h1b62, 16'h291e,
// 16'h3603, 16'h41d3, 16'h4c4b, 16'h5537,
// 16'h5c6d, 16'h61bc, 16'h6516, 16'h6665,
// 16'h6597, 16'h62c8, 16'h5dec, 16'h5730,
// 16'h4ead, 16'h4494, 16'h3912, 16'h2c71,
// 16'h1edf, 16'h10b5, 16'h022f, 16'hf3a2,
// 16'he552, 16'hd78d, 16'hca9c, 16'hbebc,
// 16'hb432, 16'hab32, 16'ha3e3, 16'h9e7e,
// 16'h9b05, 16'h99a4, 16'h9a4d, 16'h9d0d,
// 16'ha1c6, 16'ha871, 16'hb0db, 16'hbae2,
// 16'hc653, 16'hd2e8, 16'he06f, 16'hee92,
// 16'hfd17, 16'h0ba3, 16'h19fc, 16'h27c5,
// 16'h34c6, 16'h40b2, 16'h4b51, 16'h5465,
// 16'h5bc9, 16'h614c, 16'h64d7, 16'h665b,
// 16'h65c4, 16'h6327, 16'h5e7f, 16'h57f1,
// 16'h4f9b, 16'h45a5, 16'h3a4a, 16'h2dbd,
// 16'h2045, 16'h1223, 16'h03a7, 16'hf512,
// 16'he6bd, 16'hd8e5, 16'hcbdb, 16'hbfe0,
// 16'hb52d, 16'hac05, 16'ha48c, 16'h9eee,
// 16'h9b4a, 16'h99ac, 16'h9a26, 16'h9caf,
// 16'ha136, 16'ha7b2, 16'hafef, 16'hb9d1,
// 16'hc521, 16'hd197, 16'hdf0f, 16'hed21,
// 16'hfba2, 16'h0a32, 16'h188f, 16'h266d,
// 16'h3385, 16'h3f8d, 16'h4a54, 16'h538e,
// 16'h5b23, 16'h60d1, 16'h6498, 16'h6648,
// 16'h65ee, 16'h6381, 16'h5f0a, 16'h58b2,
// 16'h5080, 16'h46b9, 16'h3b78, 16'h2f0d,
// 16'h21a4, 16'h1394, 16'h051b, 16'hf687,
// 16'he827, 16'hda3f, 16'hcd1e, 16'hc104,
// 16'hb630, 16'hacdc, 16'ha535, 16'h9f69,
// 16'h9b8f, 16'h99be, 16'h9a04, 16'h9c52,
// 16'ha0b0, 16'ha6f4, 16'haf0a, 16'hb8c3,
// 16'hc3ee, 16'hd050, 16'hdda9, 16'hebb8,
// 16'hfa27, 16'h08c2, 16'h1722, 16'h2513,
// 16'h3240, 16'h3e68, 16'h494e, 16'h52b7,
// 16'h5a74, 16'h6058, 16'h644c, 16'h6637,
// 16'h660d, 16'h63d6, 16'h5f97, 16'h5964,
// 16'h516b, 16'h47c0, 16'h3caa, 16'h3055,
// 16'h2306, 16'h1501, 16'h068f, 16'hf7fd,
// 16'he991, 16'hdb9c, 16'hce65, 16'hc228,
// 16'hb73a, 16'hadb2, 16'ha5eb, 16'h9fe1,
// 16'h9bdf, 16'h99d2, 16'h99e6, 16'h9c20,
// 16'ha028, 16'ha63f, 16'hae26, 16'hb7bb,
// 16'hc2bf, 16'hcf08, 16'hdc4b, 16'hea47,
// 16'hf8b7, 16'h074a, 16'h15b7, 16'h23b7,
// 16'h30f7, 16'h3d41, 16'h4846, 16'h51d8,
// 16'h59c4, 16'h5fd5, 16'h6401, 16'h661a,
// 16'h662d, 16'h6424, 16'h601b, 16'h5a18,
// 16'h524b, 16'h48c9, 16'h3dd6, 16'h319c,
// 16'h2463, 16'h1670, 16'h0802, 16'hf973,
// 16'heafc, 16'hdcfc, 16'hcfaa, 16'hc358,
// 16'hb83d, 16'hae97, 16'ha69b, 16'ha069,
// 16'h9c2b, 16'h99f2, 16'h99c9, 16'h9bb5,
// 16'h9fa6, 16'ha58e, 16'had47, 16'hb6b5,
// 16'hc196, 16'hcdc0, 16'hdaee, 16'he8dc,
// 16'hf740, 16'h05d8, 16'h1448, 16'h2257,
// 16'h2fb1, 16'h3c10, 16'h473e, 16'h50f6,
// 16'h590b, 16'h5f52, 16'h63ad, 16'h65fb,
// 16'h6645, 16'h646e, 16'h6099, 16'h5ac9,
// 16'h5326, 16'h49ce, 16'h3eff, 16'h32e0,
// 16'h25c0, 16'h17dc, 16'h0976, 16'hfae7,
// 16'hec6c, 16'hde5b, 16'hd0f4, 16'hc487,
// 16'hb949, 16'haf7d, 16'ha752, 16'ha0f2,
// 16'h9c80, 16'h9a15, 16'h99b3, 16'h9b6d,
// 16'h9f2a, 16'ha4e0, 16'hac70, 16'hb5b0,
// 16'hc06e, 16'hcc7f, 16'hd98f, 16'he774,
// 16'hf5cc, 16'h0461, 16'h12db, 16'h20f5,
// 16'h2e66, 16'h3ae0, 16'h4630, 16'h500f,
// 16'h584f, 16'h5eca, 16'h6350, 16'h65dd,
// 16'h6650, 16'h64b9, 16'h610f, 16'h5b77,
// 16'h53fa, 16'h4ad2, 16'h4021, 16'h3425,
// 16'h271b, 16'h1944, 16'h0aeb, 16'hfc5d,
// 16'hedd9, 16'hdfbe, 16'hd242, 16'hc5b5,
// 16'hba5e, 16'hb061, 16'ha812, 16'ha17e,
// 16'h9cdd, 16'h9a38, 16'h99a8, 16'h9b27,
// 16'h9eb5, 16'ha437, 16'hab9b, 16'hb4af,
// 16'hbf4e, 16'hcb3b, 16'hd839, 16'he606,
// 16'hf45c, 16'h02e9, 16'h116f, 16'h1f90,
// 16'h2d19, 16'h39ac, 16'h451f, 16'h4f24,
// 16'h5790, 16'h5e3a, 16'h62f1, 16'h65b6,
// 16'h665b, 16'h64fa, 16'h6185, 16'h5c19,
// 16'h54d1, 16'h4bcd, 16'h4144, 16'h3564,
// 16'h2874, 16'h1aac, 16'h0c61, 16'hfdce,
// 16'hef4e, 16'he11c, 16'hd395, 16'hc6ea,
// 16'hbb6e, 16'hb152, 16'ha8d0, 16'ha213,
// 16'h9d3c, 16'h9a64, 16'h999e, 16'h9ae9,
// 16'h9e43, 16'ha394, 16'haaca, 16'hb3b2,
// 16'hbe31, 16'hc9f9, 16'hd6e5, 16'he49c,
// 16'hf2e9, 16'h0174, 16'h0ffd, 16'h1e2e,
// 16'h2bc7, 16'h3877, 16'h4409, 16'h4e34,
// 16'h56ce, 16'h5da3, 16'h6291, 16'h6586,
// 16'h6661, 16'h6538, 16'h61f1, 16'h5cbe,
// 16'h559c, 16'h4cc9, 16'h4261, 16'h36a1,
// 16'h29ca, 16'h1c15, 16'h0dd1, 16'hff47,
// 16'hf0bb, 16'he285, 16'hd4e3, 16'hc824,
// 16'hbc84, 16'hb244, 16'ha996, 16'ha2aa,
// 16'h9da0, 16'h9a97, 16'h9999, 16'h9ab1,
// 16'h9dd5, 16'ha2f7, 16'ha9fb, 16'hb2be,
// 16'hbd12, 16'hc8be, 16'hd590, 16'he335,
// 16'hf176, 16'h2001, 16'h0e89, 16'h1ccb,
// 16'h2a71, 16'h3741, 16'h42ee, 16'h4d43,
// 16'h5605, 16'h5d07, 16'h622f, 16'h654a,
// 16'h666c, 16'h6565, 16'h6262, 16'h5d55,
// 16'h566b, 16'h4dbb, 16'h437d, 16'h37dc,
// 16'h2b1c, 16'h1d7e, 16'h0f40, 16'h20be,
// 16'hf22d, 16'he3eb, 16'hd637, 16'hc95e,
// 16'hbd9e, 16'hb33a, 16'haa62, 16'ha343,
// 16'h9e0e, 16'h9ac9, 16'h999e, 16'h9a7b,
// 16'h9d6f, 16'ha25c, 16'ha933, 16'hb1cb,
// 16'hbbf9, 16'hc786, 16'hd43b, 16'he1d1,
// 16'hf003, 16'hfe8e, 16'h0d15, 16'h1b65,
// 16'h291b, 16'h3605, 16'h41d2, 16'h4c4c,
// 16'h5537, 16'h5c6b, 16'h61be, 16'h6516,
// 16'h6663, 16'h6599, 16'h62c7, 16'h5deb,
// 16'h5732, 16'h4eac, 16'h4493, 16'h3914,
// 16'h2c6f, 16'h1edf, 16'h10b6, 16'h022f,
// 16'hf3a1, 16'he553, 16'hd78d, 16'hca9b,
// 16'hbebe, 16'hb430, 16'hab33, 16'ha3e3,
// 16'h9e7e, 16'h9b06, 16'h99a2, 16'h9a4f,
// 16'h9d0a, 16'ha1c9, 16'ha86f, 16'hb0dc,
// 16'hbae2, 16'hc652, 16'hd2e9, 16'he06e,
// 16'hee93, 16'hfd15, 16'h0ba7, 16'h19f7,
// 16'h27ca, 16'h34c1, 16'h40b6, 16'h4b4e,
// 16'h5468, 16'h5bc6, 16'h614d, 16'h64d8,
// 16'h6658, 16'h65c9, 16'h6322, 16'h5e82,
// 16'h57f0, 16'h4f9b, 16'h45a6, 16'h3a4a,
// 16'h2dbc, 16'h2045, 16'h1224, 16'h03a5,
// 16'hf515, 16'he6bb, 16'hd8e5, 16'hcbdd,
// 16'hbfdc, 16'hb531, 16'hac03, 16'ha48c,
// 16'h9ef0, 16'h9b47, 16'h99ae, 16'h9a27,
// 16'h9cab, 16'ha13c, 16'ha7ac, 16'haff3,
// 16'hb9d0, 16'hc51f, 16'hd19b, 16'hdf0c,
// 16'hed22, 16'hfba1, 16'h0a32, 16'h1890,
// 16'h266c, 16'h3386, 16'h3f8c, 16'h4a54,
// 16'h538f, 16'h5b21, 16'h60d4, 16'h6496,
// 16'h6648, 16'h65f0, 16'h637d, 16'h5f10,
// 16'h58ac, 16'h5085, 16'h46b5, 16'h3b7b,
// 16'h2f0a, 16'h21a7, 16'h1392, 16'h051c,
// 16'hf686, 16'he828, 16'hda3f, 16'hcd1d,
// 16'hc106, 16'hb62c, 16'hace1, 16'ha531,
// 16'h9f6c, 16'h9b8d, 16'h99c0, 16'h9a20,
// 16'h9c57, 16'ha0ac, 16'ha6f6, 16'haf0a,
// 16'hb8c1, 16'hc3f0, 16'hd04f, 16'hddab,
// 16'hebb4, 16'hfa2c, 16'h08bd, 16'h1726,
// 16'h2511, 16'h3240, 16'h3e69, 16'h494e,
// 16'h52b7, 16'h5a73, 16'h6058, 16'h644e,
// 16'h6634, 16'h6611, 16'h63d2, 16'h5f9a,
// 16'h5963, 16'h516b, 16'h47c0, 16'h3caa,
// 16'h3055, 16'h2306, 16'h1520, 16'h0692,
// 16'hf7f9, 16'he994, 16'hdb9b, 16'hce63,
// 16'hc22d, 16'hb733, 16'hadba, 16'ha5e2,
// 16'h9feb, 16'h9bd7, 16'h99d7, 16'h99e3,
// 16'h9c01, 16'ha029, 16'ha63e, 16'hae28,
// 16'hb7b8, 16'hc2c1, 16'hcf08, 16'hdc49,
// 16'hea4a, 16'hf8b4, 16'h074c, 16'h15b7,
// 16'h23b5, 16'h30f9, 16'h3d3f, 16'h4847,
// 16'h51db, 16'h59bd, 16'h5fdd, 16'h63fa,
// 16'h6620, 16'h6629, 16'h6425, 16'h601b,
// 16'h5a19, 16'h524a, 16'h48ca, 16'h3dd5,
// 16'h319b, 16'h2467, 16'h166b, 16'h0807,
// 16'hf96e, 16'heb20, 16'hdcfa, 16'hcfab,
// 16'hc357, 16'hb83d, 16'hae99, 16'ha698,
// 16'ha06b, 16'h9c2b, 16'h99f0, 16'h99cc,
// 16'h9bb1, 16'h9fa9, 16'ha58d, 16'had48,
// 16'hb6b4, 16'hc194, 16'hcdc4, 16'hdaea,
// 16'he8e0, 16'hf73e, 16'h05d7, 16'h144a,
// 16'h2256, 16'h2fb1, 16'h3c10, 16'h473f,
// 16'h50f4, 16'h590d, 16'h5f51, 16'h63ac,
// 16'h65fe, 16'h6641, 16'h6471, 16'h6098,
// 16'h5ac9, 16'h5326, 16'h49cf, 16'h3efc,
// 16'h32e3, 16'h25bf, 16'h17db, 16'h0978,
// 16'hfae5, 16'hec6d, 16'hde5a, 16'hd0f6,
// 16'hc484, 16'hb94c, 16'haf7b, 16'ha752,
// 16'ha0f4, 16'h9c7d, 16'h9a17, 16'h99b2,
// 16'h9b6e, 16'h9f2a, 16'ha4e0, 16'hac6f,
// 16'hb5af, 16'hc071, 16'hcc7c, 16'hd993,
// 16'he770, 16'hf5cd, 16'h0462, 16'h12d9,
// 16'h20f9, 16'h2e60, 16'h3ae6, 16'h462b,
// 16'h5013, 16'h584e, 16'h5ec7, 16'h6354,
// 16'h65d9, 16'h6655, 16'h64b4, 16'h6114,
// 16'h5b72, 16'h53fd, 16'h4ad2, 16'h4020,
// 16'h3426, 16'h271a, 16'h1945, 16'h0aea,
// 16'hfc5d, 16'hedda, 16'hdfbd, 16'hd242,
// 16'hc5b7, 16'hba59, 16'hb067, 16'ha80d,
// 16'ha181, 16'h9cdb, 16'h9a39, 16'h99a8,
// 16'h9b26, 16'h9eb6, 16'ha436, 16'hab9c,
// 16'hb4ae, 16'hbf4f, 16'hcb39, 16'hd83b,
// 16'he605, 16'hf45c, 16'h02ea, 16'h116c,
// 16'h1f94, 16'h2d14, 16'h39b2, 16'h4519,
// 16'h4f29, 16'h578c, 16'h5e3c, 16'h62f2,
// 16'h65b4, 16'h665c, 16'h64fa, 16'h6183,
// 16'h5c1d, 16'h54cd, 16'h4bd0, 16'h4142,
// 16'h3564, 16'h2875, 16'h1aab, 16'h0c62,
// 16'hfdcd, 16'hef4e, 16'he11d, 16'hd394,
// 16'hc6ea, 16'hbb6e, 16'hb153, 16'ha8cf,
// 16'ha213, 16'h9d3c, 16'h9a63, 16'h99a1,
// 16'h9ae6, 16'h9e45, 16'ha394, 16'haac8,
// 16'hb3b6, 16'hbe2c, 16'hc9fe, 16'hd6e0,
// 16'he4a0, 16'hf2e7, 16'h0175, 16'h0ffd,
// 16'h1e2d, 16'h2bc6, 16'h387a, 16'h4406,
// 16'h4e38, 16'h56ca, 16'h5da5, 16'h6291,
// 16'h6585, 16'h6663, 16'h6535, 16'h61f4,
// 16'h5cbb, 16'h559f, 16'h4cc7, 16'h4260,
// 16'h36a4, 16'h29c7, 16'h1c17, 16'h0dcf,
// 16'hff49, 16'hf0b8, 16'he28a, 16'hd4de,
// 16'hc827, 16'hbc82, 16'hb244, 16'ha999,
// 16'ha2a6, 16'h9da4, 16'h9a93, 16'h999c,
// 16'h9ab0, 16'h9dd5, 16'ha2f6, 16'ha9fd,
// 16'hb2bc, 16'hbd13, 16'hc8bf, 16'hd58d,
// 16'he338, 16'hf174, 16'h2002, 16'h0e88,
// 16'h1ccc, 16'h2a6f, 16'h3744, 16'h42eb,
// 16'h4d46, 16'h5602, 16'h5d09, 16'h622d,
// 16'h654c, 16'h666b, 16'h6565, 16'h6263,
// 16'h5d54, 16'h566c, 16'h4dba, 16'h437d,
// 16'h37dd, 16'h2b1b, 16'h1d7e, 16'h0f42,
// 16'h20ba, 16'hf231, 16'he3e8, 16'hd639,
// 16'hc95d, 16'hbd9e, 16'hb33c, 16'haa5e,
// 16'ha348, 16'h9e09, 16'h9acd, 16'h999c,
// 16'h9a7c, 16'h9d6e, 16'ha25c, 16'ha935,
// 16'hb1c8, 16'hbbfb, 16'hc785, 16'hd43b,
// 16'he1d2, 16'hf003, 16'hfe8c, 16'h0d18,
// 16'h1b61, 16'h291f, 16'h3603, 16'h41d2,
// 16'h4c4d, 16'h5535, 16'h5c6e, 16'h61bc,
// 16'h6517, 16'h6662, 16'h659b, 16'h62c5,
// 16'h5dee, 16'h572f, 16'h4eae, 16'h4492,
// 16'h3915, 16'h2c6e, 16'h1ee1, 16'h10b4,
// 16'h0231, 16'hf39f, 16'he555, 16'hd78a,
// 16'hca9f, 16'hbeba, 16'hb434, 16'hab2f,
// 16'ha3e6, 16'h9e7c, 16'h9b06, 16'h99a3,
// 16'h9a4e, 16'h9d0a, 16'ha1ca, 16'ha86e,
// 16'hb0dc, 16'hbae3, 16'hc650, 16'hd2eb,
// 16'he06d, 16'hee94, 16'hfd15, 16'h0ba5,
// 16'h19f9, 16'h27c8, 16'h34c4, 16'h40b4,
// 16'h4b4e, 16'h5468, 16'h5bc7, 16'h614c,
// 16'h64d9, 16'h6658, 16'h65c6, 16'h6327,
// 16'h5e7e, 16'h57f2, 16'h4f9a, 16'h45a7,
// 16'h3a47, 16'h2dc1, 16'h2040, 16'h1228,
// 16'h03a3, 16'hf515, 16'he6bb, 16'hd8e7,
// 16'hcbd8, 16'hbfe2, 16'hb52d, 16'hac05,
// 16'ha48b, 16'h9eee, 16'h9b4a, 16'h99ae,
// 16'h9a25, 16'h9cad, 16'ha139, 16'ha7af,
// 16'haff2, 16'hb9cf, 16'hc521, 16'hd198,
// 16'hdf0f, 16'hed21, 16'hfba1, 16'h0a32,
// 16'h188f, 16'h266e, 16'h3384, 16'h3f8f,
// 16'h4a51, 16'h5390, 16'h5b21, 16'h60d4,
// 16'h6496, 16'h6649, 16'h65ee, 16'h637f,
// 16'h5f0e, 16'h58ae, 16'h5083, 16'h46b7,
// 16'h3b79, 16'h2f0d, 16'h21a3, 16'h1396,
// 16'h0517, 16'hf68c, 16'he822, 16'hda44,
// 16'hcd1a, 16'hc106, 16'hb62f, 16'hacdc,
// 16'ha537, 16'h9f67, 16'h9b90, 16'h99be,
// 16'h9a03, 16'h9c54, 16'ha0ae, 16'ha6f6,
// 16'haf08, 16'hb8c5, 16'hc3ec, 16'hd052,
// 16'hdda8, 16'hebb8, 16'hfa28, 16'h08c1,
// 16'h1722, 16'h2514, 16'h323f, 16'h3e69,
// 16'h494e, 16'h52b6, 16'h5a75, 16'h6057,
// 16'h644e, 16'h6635, 16'h660e, 16'h63d7,
// 16'h5f94, 16'h5969, 16'h5165, 16'h47c6,
// 16'h3ca5, 16'h3059, 16'h2303, 16'h1502,
// 16'h0691, 16'hf7fa, 16'he992, 16'hdb9d,
// 16'hce63, 16'hc22b, 16'hb736, 16'hadb6,
// 16'ha5e7, 16'h9fe6, 16'h9bdb, 16'h99d4,
// 16'h99e5, 16'h9c20, 16'ha02a, 16'ha63c,
// 16'hae2a, 16'hb7b7, 16'hc2c2, 16'hcf07,
// 16'hdc49, 16'hea4a, 16'hf8b5, 16'h074b,
// 16'h15b7, 16'h23b5, 16'h30f9, 16'h3d3f,
// 16'h4849, 16'h51d6, 16'h59c4, 16'h5fd4,
// 16'h6403, 16'h661a, 16'h662c, 16'h6424,
// 16'h601b, 16'h5a19, 16'h524a, 16'h48c9,
// 16'h3dd6, 16'h319c, 16'h2465, 16'h166d,
// 16'h0805, 16'hf970, 16'heaff, 16'hdcfa,
// 16'hcfab, 16'hc358, 16'hb83d, 16'hae98,
// 16'ha699, 16'ha06a, 16'h9c2c, 16'h99f0,
// 16'h99cc, 16'h9bb1, 16'h9faa, 16'ha58a,
// 16'had4c, 16'hb6b0, 16'hc199, 16'hcdbe,
// 16'hdaf0, 16'he8da, 16'hf743, 16'h05d5,
// 16'h1448, 16'h225a, 16'h2fac, 16'h3c16,
// 16'h473b, 16'h50f5, 16'h590d, 16'h5f51,
// 16'h63ac, 16'h65fe, 16'h6642, 16'h646f,
// 16'h609a, 16'h5ac7, 16'h5328, 16'h49cc,
// 16'h3f20, 16'h32e0, 16'h25c0, 16'h17db,
// 16'h0977, 16'hfae7, 16'hec6c, 16'hde5a,
// 16'hd0f6, 16'hc485, 16'hb94a, 16'haf7d,
// 16'ha751, 16'ha0f5, 16'h9c7c, 16'h9a18,
// 16'h99b1, 16'h9b6f, 16'h9f29, 16'ha4e1,
// 16'hac6f, 16'hb5b0, 16'hc06f, 16'hcc7e,
// 16'hd991, 16'he772, 16'hf5cd, 16'h0460,
// 16'h12db, 16'h20f7, 16'h2e63, 16'h3ae3,
// 16'h462d, 16'h5011, 16'h584f, 16'h5ec9,
// 16'h6351, 16'h65db, 16'h6653, 16'h64b6,
// 16'h6113, 16'h5b72, 16'h53fd, 16'h4ad1,
// 16'h4021, 16'h3425, 16'h271a, 16'h1945,
// 16'h0aeb, 16'hfc5c, 16'hedda, 16'hdfbd,
// 16'hd243, 16'hc5b6, 16'hba5b, 16'hb064,
// 16'ha810, 16'ha180, 16'h9cdb, 16'h9a3a,
// 16'h99a6, 16'h9b29, 16'h9eb2, 16'ha43b,
// 16'hab97, 16'hb4b3, 16'hbf4a, 16'hcb3d,
// 16'hd838, 16'he608, 16'hf45a, 16'h02eb,
// 16'h116b, 16'h1f95, 16'h2d13, 16'h39b2,
// 16'h451b, 16'h4f26, 16'h578f, 16'h5e39,
// 16'h62f4, 16'h65b3, 16'h665d, 16'h64f8,
// 16'h6186, 16'h5c1a, 16'h54d0, 16'h4bcc,
// 16'h4146, 16'h3562, 16'h2874, 16'h1aae,
// 16'h0c5e, 16'hfdd1, 16'hef4b, 16'he11f,
// 16'hd392, 16'hc6ec, 16'hbb6d, 16'hb153,
// 16'ha8d0, 16'ha213, 16'h9d3a, 16'h9a66,
// 16'h999d, 16'h9aeb, 16'h9e40, 16'ha398,
// 16'haac5, 16'hb3b7, 16'hbe2d, 16'hc9fc,
// 16'hd6e2, 16'he49f, 16'hf2e7, 16'h0175,
// 16'h0ffd, 16'h1e2e, 16'h2bc6, 16'h3879,
// 16'h4407, 16'h4e35, 16'h56ce, 16'h5da2,
// 16'h6295, 16'h6580, 16'h6667, 16'h6531,
// 16'h61f8, 16'h5cb9, 16'h55a0, 16'h4cc6,
// 16'h4261, 16'h36a4, 16'h29c6, 16'h1c18,
// 16'h0dd0, 16'hff45, 16'hf0bf, 16'he280,
// 16'hd4e8, 16'hc81f, 16'hbc88, 16'hb241,
// 16'ha999, 16'ha2a7, 16'h9da3, 16'h9a93,
// 16'h999d, 16'h9aaf, 16'h9dd6, 16'ha2f5,
// 16'ha9fe, 16'hb2ba, 16'hbd16, 16'hc8bc,
// 16'hd590, 16'he335, 16'hf178, 16'hfffc,
// 16'h0e8f, 16'h1cc6, 16'h2a74, 16'h3741,
// 16'h42ec, 16'h4d45, 16'h5602, 16'h5d0c,
// 16'h6228, 16'h6553, 16'h6663, 16'h656b,
// 16'h6261, 16'h5d53, 16'h566e, 16'h4db8,
// 16'h437f, 16'h37da, 16'h2b1f, 16'h1d7a,
// 16'h0f44, 16'h20bb, 16'hf22e, 16'he3eb,
// 16'hd637, 16'hc95d, 16'hbda0, 16'hb339,
// 16'haa61, 16'ha345, 16'h9e0b, 16'h9acc,
// 16'h999d, 16'h9a7b, 16'h9d6f, 16'ha25b,
// 16'ha935, 16'hb1c9, 16'hbbfb, 16'hc785,
// 16'hd43a, 16'he1d3, 16'hf001, 16'hfe90,
// 16'h0d13, 16'h1b65, 16'h291c, 16'h3605,
// 16'h41d1, 16'h4c4d, 16'h5536, 16'h5c6c,
// 16'h61bd, 16'h6517, 16'h6662, 16'h659b,
// 16'h62c5, 16'h5ded, 16'h5730, 16'h4ead,
// 16'h4494, 16'h3912, 16'h2c71, 16'h1ede,
// 16'h10b7, 16'h022e, 16'hf3a2, 16'he552,
// 16'hd78d, 16'hca9c, 16'hbebc, 16'hb433,
// 16'hab30, 16'ha3e7, 16'h9e79, 16'h9b08,
// 16'h99a3, 16'h9a4d, 16'h9d0d, 16'ha1c7,
// 16'ha86e, 16'hb0de, 16'hbae1, 16'hc652,
// 16'hd2ea, 16'he06d, 16'hee93, 16'hfd17,
// 16'h0ba4, 16'h19fa, 16'h27c7, 16'h34c4,
// 16'h40b4, 16'h4b4f, 16'h5467, 16'h5bc7,
// 16'h614d, 16'h64d8, 16'h6658, 16'h65c8,
// 16'h6323, 16'h5e82, 16'h57f0, 16'h4f9b,
// 16'h45a6, 16'h3a49, 16'h2dbd, 16'h2045,
// 16'h1223, 16'h03a7, 16'hf513, 16'he6bc,
// 16'hd8e5, 16'hcbdc, 16'hbfde, 16'hb530,
// 16'hac03, 16'ha48c, 16'h9eef, 16'h9b49,
// 16'h99ae, 16'h9a24, 16'h9caf, 16'ha137,
// 16'ha7b2, 16'hafed, 16'hb9d6, 16'hc519,
// 16'hd1a0, 16'hdf08, 16'hed25, 16'hfba1,
// 16'h0a30, 16'h1891, 16'h266d, 16'h3384,
// 16'h3f90, 16'h4a4f, 16'h5393, 16'h5b1e,
// 16'h60d6, 16'h6494, 16'h664b, 16'h65ed,
// 16'h6380, 16'h5f0c, 16'h58b0, 16'h5081,
// 16'h46b9, 16'h3b78, 16'h2f0c, 16'h21a5,
// 16'h1394, 16'h0519, 16'hf68a, 16'he824,
// 16'hda42, 16'hcd1c, 16'hc105, 16'hb62f,
// 16'hacdd, 16'ha535, 16'h9f68, 16'h9b90,
// 16'h99bf, 16'h9a01, 16'h9c56, 16'ha0ac,
// 16'ha6f6, 16'haf0b, 16'hb8c1, 16'hc3f0,
// 16'hd04e, 16'hddac, 16'hebb4, 16'hfa2c,
// 16'h08be, 16'h1724, 16'h2512, 16'h3241,
// 16'h3e66, 16'h4953, 16'h52b1, 16'h5a78,
// 16'h6055, 16'h644f, 16'h6634, 16'h6610,
// 16'h63d5, 16'h5f95, 16'h5968, 16'h5167,
// 16'h47c3, 16'h3ca9, 16'h3055, 16'h2305,
// 16'h1503, 16'h068e, 16'hf7fd, 16'he991,
// 16'hdb9d, 16'hce62, 16'hc22c, 16'hb735,
// 16'hadb8, 16'ha5e5, 16'h9fe7, 16'h9bda,
// 16'h99d6, 16'h99e3, 16'h9c01, 16'ha02a,
// 16'ha63c, 16'hae2a, 16'hb7b7, 16'hc2c2,
// 16'hcf06, 16'hdc4b, 16'hea49, 16'hf8b5,
// 16'h074c, 16'h15b4, 16'h23b9, 16'h30f6,
// 16'h3d42, 16'h4845, 16'h51da, 16'h59c0,
// 16'h5fda, 16'h63fc, 16'h661f, 16'h6629,
// 16'h6426, 16'h601a, 16'h5a1a, 16'h5249,
// 16'h48ca, 16'h3dd5, 16'h319d, 16'h2464,
// 16'h166e, 16'h0804, 16'hf970, 16'heaff,
// 16'hdcfb, 16'hcfaa, 16'hc357, 16'hb83f,
// 16'hae95, 16'ha69d, 16'ha067, 16'h9c2d,
// 16'h99f0, 16'h99cb, 16'h9bb3, 16'h9fa8,
// 16'ha58c, 16'had4a, 16'hb6b2, 16'hc196,
// 16'hcdc3, 16'hdaea, 16'he8df, 16'hf740,
// 16'h05d6, 16'h144b, 16'h2254, 16'h2fb2,
// 16'h3c10, 16'h473f, 16'h50f6, 16'h5909,
// 16'h5f56, 16'h63a6, 16'h6604, 16'h663c,
// 16'h6475, 16'h6095, 16'h5acc, 16'h5322,
// 16'h49d3, 16'h3ef9, 16'h32e6, 16'h25bd,
// 16'h17db, 16'h0978, 16'hfae7, 16'hec6a,
// 16'hde5e, 16'hd0f0, 16'hc48b, 16'hb946,
// 16'haf80, 16'ha750, 16'ha0f2, 16'h9c82,
// 16'h9a12, 16'h99b6, 16'h9b6b, 16'h9f2b,
// 16'ha4e0, 16'hac71, 16'hb5ad, 16'hc071,
// 16'hcc7c, 16'hd993, 16'he770, 16'hf5cf,
// 16'h045f, 16'h12db, 16'h20f8, 16'h2e60,
// 16'h3ae7, 16'h462a, 16'h5014, 16'h584c,
// 16'h5ecb, 16'h634f, 16'h65de, 16'h6650,
// 16'h64b9, 16'h6110, 16'h5b75, 16'h53fb,
// 16'h4ad3, 16'h401f, 16'h3427, 16'h2719,
// 16'h1945, 16'h0aec, 16'hfc5b, 16'heddb,
// 16'hdfbc, 16'hd243, 16'hc5b5, 16'hba5d,
// 16'hb063, 16'ha810, 16'ha17f, 16'h9cdb,
// 16'h9a3b, 16'h99a6, 16'h9b28, 16'h9eb4,
// 16'ha438, 16'hab9a, 16'hb4b0, 16'hbf4d,
// 16'hcb3b, 16'hd83a, 16'he606, 16'hf45b,
// 16'h02e9, 16'h116f, 16'h1f8f, 16'h2d1b,
// 16'h39aa, 16'h4521, 16'h4f22, 16'h5792,
// 16'h5e37, 16'h62f6, 16'h65b0, 16'h6660,
// 16'h64f7, 16'h6186, 16'h5c1a, 16'h54cf,
// 16'h4bcf, 16'h4142, 16'h3566, 16'h2871,
// 16'h1ab0, 16'h0c5d, 16'hfdd1, 16'hef4c,
// 16'he11e, 16'hd393, 16'hc6eb, 16'hbb6d,
// 16'hb154, 16'ha8ce, 16'ha215, 16'h9d39,
// 16'h9a66, 16'h999e, 16'h9ae9, 16'h9e43,
// 16'ha394, 16'haaca, 16'hb3b3, 16'hbe2f,
// 16'hc9fb, 16'hd6e3, 16'he49e, 16'hf2e8,
// 16'h0175, 16'h0ffc, 16'h1e2e, 16'h2bc7,
// 16'h3877, 16'h440a, 16'h4e33, 16'h56cf,
// 16'h5da1, 16'h6294, 16'h6582, 16'h6666,
// 16'h6533, 16'h61f5, 16'h5cbb, 16'h559e,
// 16'h4cc8, 16'h4261, 16'h36a1, 16'h29cb,
// 16'h1c13, 16'h0dd3, 16'hff44, 16'hf0bf,
// 16'he281, 16'hd4e8, 16'hc81e, 16'hbc89,
// 16'hb240, 16'ha99a, 16'ha2a7, 16'h9da2,
// 16'h9a96, 16'h9998, 16'h9ab4, 16'h9dd2,
// 16'ha2f8, 16'ha9fc, 16'hb2bc, 16'hbd13,
// 16'hc8bf, 16'hd58e, 16'he337, 16'hf175,
// 16'h2020, 16'h0e8b, 16'h1cc9, 16'h2a72,
// 16'h3741, 16'h42ee, 16'h4d42, 16'h5606,
// 16'h5d07, 16'h622d, 16'h654e, 16'h6667,
// 16'h656a, 16'h625f, 16'h5d57, 16'h5668,
// 16'h4dbf, 16'h4378, 16'h37e1, 16'h2b18,
// 16'h1d7f, 16'h0f42, 16'h20ba, 16'hf230,
// 16'he3ea, 16'hd636, 16'hc95f, 16'hbd9f,
// 16'hb338, 16'haa63, 16'ha343, 16'h9e0d,
// 16'h9acb, 16'h999d, 16'h9a7a, 16'h9d70,
// 16'ha25c, 16'ha933, 16'hb1cb, 16'hbbf7,
// 16'hc789, 16'hd439, 16'he1d3, 16'hf002,
// 16'hfe8c, 16'h0d18, 16'h1b62, 16'h291e,
// 16'h3603, 16'h41d4, 16'h4c49, 16'h553a,
// 16'h5c69, 16'h61bf, 16'h6516, 16'h6662,
// 16'h659c, 16'h62c2, 16'h5df2, 16'h572a,
// 16'h4eb3, 16'h448f, 16'h3915, 16'h2c70,
// 16'h1ede, 16'h10b7, 16'h022e, 16'hf3a3,
// 16'he550, 16'hd790, 16'hca99, 16'hbebe,
// 16'hb432, 16'hab30, 16'ha3e7, 16'h9e7a,
// 16'h9b08, 16'h99a1, 16'h9a50, 16'h9d09,
// 16'ha1cb, 16'ha86d, 16'hb0dd, 16'hbae2,
// 16'hc651, 16'hd2eb, 16'he06c, 16'hee96,
// 16'hfd12, 16'h0ba8, 16'h19f8, 16'h27c7,
// 16'h34c6, 16'h40b2, 16'h4b4f, 16'h5469,
// 16'h5bc4, 16'h614f, 16'h64d7, 16'h6659,
// 16'h65c8, 16'h6322, 16'h5e82, 16'h57f0,
// 16'h4f9c, 16'h45a5, 16'h3a4a, 16'h2dbc,
// 16'h2046, 16'h1223, 16'h03a6, 16'hf514,
// 16'he6bb, 16'hd8e7, 16'hcbda, 16'hbfdf,
// 16'hb52f, 16'hac03, 16'ha48e, 16'h9eec,
// 16'h9b4b, 16'h99ac, 16'h9a27, 16'h9cac,
// 16'ha13a, 16'ha7ae, 16'haff1, 16'hb9d3,
// 16'hc51b, 16'hd19f, 16'hdf08, 16'hed26,
// 16'hfb9f, 16'h0a32, 16'h1890, 16'h266d,
// 16'h3384, 16'h3f90, 16'h4a50, 16'h5391,
// 16'h5b20, 16'h60d5, 16'h6495, 16'h664a,
// 16'h65ed, 16'h6380, 16'h5f0d, 16'h58b0,
// 16'h5081, 16'h46b8, 16'h3b7a, 16'h2f09,
// 16'h21a9, 16'h1390, 16'h051d, 16'hf687,
// 16'he825, 16'hda41, 16'hcd1d, 16'hc104,
// 16'hb630, 16'hacdc, 16'ha535, 16'h9f69,
// 16'h9b8f, 16'h99be, 16'h9a04, 16'h9c52,
// 16'ha0b0, 16'ha6f3, 16'haf0b, 16'hb8c3,
// 16'hc3ee, 16'hd050, 16'hdda9, 16'hebb8,
// 16'hfa27, 16'h08c3, 16'h171f, 16'h2517,
// 16'h323d, 16'h3e6a, 16'h494d, 16'h52b8,
// 16'h5a71, 16'h605c, 16'h6449, 16'h6639,
// 16'h660c, 16'h63d7, 16'h5f95, 16'h5968,
// 16'h5166, 16'h47c4, 16'h3ca8, 16'h3056,
// 16'h2305, 16'h1501, 16'h0690, 16'hf7fb,
// 16'he994, 16'hdb99, 16'hce66, 16'hc22a,
// 16'hb734, 16'hadba, 16'ha5e3, 16'h9fe9,
// 16'h9bd9, 16'h99d6, 16'h99e2, 16'h9c03,
// 16'ha027, 16'ha640, 16'hae26, 16'hb7ba,
// 16'hc2c0, 16'hcf08, 16'hdc4a, 16'hea49,
// 16'hf8b4, 16'h074d, 16'h15b6, 16'h23b5,
// 16'h30fa, 16'h3d3d, 16'h484a, 16'h51d7,
// 16'h59c2, 16'h5fd7, 16'h63ff, 16'h661c,
// 16'h662c, 16'h6425, 16'h601a, 16'h5a19,
// 16'h5249, 16'h48cb, 16'h3dd5, 16'h319c,
// 16'h2465, 16'h166c, 16'h0807, 16'hf96d,
// 16'heb02, 16'hdcf8, 16'hcfac, 16'hc358,
// 16'hb83b, 16'hae9b, 16'ha697, 16'ha06b,
// 16'h9c2b, 16'h99f1, 16'h99ca, 16'h9bb4,
// 16'h9fa7, 16'ha58c, 16'had4b, 16'hb6b0,
// 16'hc199, 16'hcdbf, 16'hdaee, 16'he8db,
// 16'hf743, 16'h05d5, 16'h144a, 16'h2256,
// 16'h2fb0, 16'h3c12, 16'h473e, 16'h50f5,
// 16'h590c, 16'h5f51, 16'h63ac, 16'h65fe,
// 16'h6641, 16'h6472, 16'h6096, 16'h5acc,
// 16'h5322, 16'h49d3, 16'h3ef9, 16'h32e5,
// 16'h25be, 16'h17dc, 16'h0978, 16'hfae4,
// 16'hec6f, 16'hde57, 16'hd0f8, 16'hc485,
// 16'hb948, 16'haf81, 16'ha74d, 16'ha0f5,
// 16'h9c80, 16'h9a13, 16'h99b6, 16'h9b6b,
// 16'h9f2a, 16'ha4e2, 16'hac6f, 16'hb5ad,
// 16'hc075, 16'hcc76, 16'hd999, 16'he76b,
// 16'hf5d1, 16'h0460, 16'h12db, 16'h20f6,
// 16'h2e63, 16'h3ae3, 16'h462e, 16'h5011,
// 16'h584f, 16'h5ec8, 16'h6353, 16'h65da,
// 16'h6653, 16'h64b6, 16'h6113, 16'h5b73,
// 16'h53fe, 16'h4ace, 16'h4024, 16'h3424,
// 16'h271a, 16'h1946, 16'h0ae9, 16'hfc5d,
// 16'heddc, 16'hdfba, 16'hd245, 16'hc5b4,
// 16'hba5c, 16'hb065, 16'ha80f, 16'ha180,
// 16'h9cdb, 16'h9a3a, 16'h99a5, 16'h9b2b,
// 16'h9eb1, 16'ha43b, 16'hab98, 16'hb4af,
// 16'hbf50, 16'hcb38, 16'hd83c, 16'he605,
// 16'hf45a, 16'h02ed, 16'h1169, 16'h1f97,
// 16'h2d12, 16'h39b2, 16'h451b, 16'h4f25,
// 16'h5791, 16'h5e38, 16'h62f5, 16'h65b1,
// 16'h665f, 16'h64f6, 16'h6189, 16'h5c17,
// 16'h54d1, 16'h4bcf, 16'h413f, 16'h356a,
// 16'h286f, 16'h1aaf, 16'h0c60, 16'hfdcd,
// 16'hef4e, 16'he11f, 16'hd391, 16'hc6ed,
// 16'hbb6b, 16'hb154, 16'ha8d1, 16'ha211,
// 16'h9d3c, 16'h9a65, 16'h999e, 16'h9ae9,
// 16'h9e43, 16'ha393, 16'haacb, 16'hb3b3,
// 16'hbe2e, 16'hc9fc, 16'hd6e3, 16'he49c,
// 16'hf2ea, 16'h0173, 16'h0ffd, 16'h1e2f,
// 16'h2bc5, 16'h3879, 16'h4407, 16'h4e37,
// 16'h56ca, 16'h5da7, 16'h628f, 16'h6585,
// 16'h6665, 16'h6532, 16'h61f7, 16'h5cb9,
// 16'h55a0, 16'h4cc6, 16'h4262, 16'h36a1,
// 16'h29ca, 16'h1c15, 16'h0dd1, 16'hff46,
// 16'hf0bd, 16'he283, 16'hd4e4, 16'hc824,
// 16'hbc83, 16'hb245, 16'ha996, 16'ha2a9,
// 16'h9da1, 16'h9a96, 16'h999a, 16'h9ab0,
// 16'h9dd7, 16'ha2f3, 16'haa20, 16'hb2b9,
// 16'hbd16, 16'hc8bc, 16'hd590, 16'he335,
// 16'hf177, 16'hffff, 16'h0e8b, 16'h1cc9,
// 16'h2a72, 16'h3740, 16'h42f0, 16'h4d40,
// 16'h5607, 16'h5d07, 16'h622d, 16'h654e,
// 16'h6667, 16'h6569, 16'h6260, 16'h5d57,
// 16'h5669, 16'h4dbd, 16'h437a, 16'h37df,
// 16'h2b1a, 16'h1d7e, 16'h0f42, 16'h20bb,
// 16'hf22e, 16'he3eb, 16'hd637, 16'hc95e,
// 16'hbd9e, 16'hb33b, 16'haa5e, 16'ha349,
// 16'h9e08, 16'h9ace, 16'h999b, 16'h9a7c,
// 16'h9d6e, 16'ha25e, 16'ha931, 16'hb1cd,
// 16'hbbf5, 16'hc78a, 16'hd439, 16'he1d2,
// 16'hf004, 16'hfe8a, 16'h0d19, 16'h1b61,
// 16'h291f, 16'h3602, 16'h41d5, 16'h4c49,
// 16'h5539, 16'h5c6a, 16'h61be, 16'h6517,
// 16'h6662, 16'h659b, 16'h62c4, 16'h5def,
// 16'h572d, 16'h4eb0, 16'h4491, 16'h3915,
// 16'h2c6f, 16'h1edf, 16'h10b5, 16'h0230,
// 16'hf3a2, 16'he551, 16'hd790, 16'hca98,
// 16'hbebf, 16'hb432, 16'hab2f, 16'ha3e8,
// 16'h9e79, 16'h9b09, 16'h99a1, 16'h9a4e,
// 16'h9d0c, 16'ha1c8, 16'ha86e, 16'hb0de,
// 16'hbadf, 16'hc655, 16'hd2e8, 16'he06e,
// 16'hee93, 16'hfd16, 16'h0ba4, 16'h19fc,
// 16'h27c5, 16'h34c5, 16'h40b4, 16'h4b4f,
// 16'h5466, 16'h5bca, 16'h6148, 16'h64dd,
// 16'h6655, 16'h65ca, 16'h6321, 16'h5e83,
// 16'h57f0, 16'h4f9b, 16'h45a6, 16'h3a49,
// 16'h2dbc, 16'h2046, 16'h1223, 16'h03a6,
// 16'hf515, 16'he6ba, 16'hd8e6, 16'hcbdb,
// 16'hbfdf, 16'hb52f, 16'hac04, 16'ha48c,
// 16'h9eed, 16'h9b4c, 16'h99aa, 16'h9a28,
// 16'h9cad, 16'ha137, 16'ha7b2, 16'hafef,
// 16'hb9d1, 16'hc520, 16'hd19a, 16'hdf0b,
// 16'hed25, 16'hfb9e, 16'h0a35, 16'h188d,
// 16'h2670, 16'h3381, 16'h3f92, 16'h4a4f,
// 16'h5392, 16'h5b1f, 16'h60d6, 16'h6493,
// 16'h664e, 16'h65e8, 16'h6384, 16'h5f0b,
// 16'h58af, 16'h5083, 16'h46b6, 16'h3b7a,
// 16'h2f0d, 16'h21a3, 16'h1395, 16'h0519,
// 16'hf689, 16'he826, 16'hda40, 16'hcd1e,
// 16'hc102, 16'hb632, 16'hacda, 16'ha538,
// 16'h9f67, 16'h9b8f, 16'h99bf, 16'h9a01,
// 16'h9c56, 16'ha0ad, 16'ha6f6, 16'haf09,
// 16'hb8c3, 16'hc3ee, 16'hd050, 16'hddaa,
// 16'hebb6, 16'hfa2b, 16'h08be, 16'h1724,
// 16'h2511, 16'h3243, 16'h3e65, 16'h4953,
// 16'h52b1, 16'h5a78, 16'h6055, 16'h6450,
// 16'h6633, 16'h6611, 16'h63d4, 16'h5f96,
// 16'h5967, 16'h5168, 16'h47c2, 16'h3caa,
// 16'h3055, 16'h2304, 16'h1504, 16'h068c,
// 16'hf820, 16'he98e, 16'hdba0, 16'hce5f,
// 16'hc22f, 16'hb733, 16'hadb8, 16'ha5e6,
// 16'h9fe6, 16'h9bda, 16'h99d7, 16'h99e2,
// 16'h9c01, 16'ha02a, 16'ha63b, 16'hae2c,
// 16'hb7b5, 16'hc2c4, 16'hcf04, 16'hdc4c,
// 16'hea49, 16'hf8b4, 16'h074d, 16'h15b4,
// 16'h23b9, 16'h30f6, 16'h3d42, 16'h4844,
// 16'h51db, 16'h59c0, 16'h5fd9, 16'h63fe,
// 16'h661e, 16'h6629, 16'h6426, 16'h601a,
// 16'h5a19, 16'h524c, 16'h48c7, 16'h3dd8,
// 16'h319a, 16'h2466, 16'h166d, 16'h0805,
// 16'hf96f, 16'heb01, 16'hdcf8, 16'hcfad,
// 16'hc356, 16'hb83d, 16'hae99, 16'ha699,
// 16'ha06a, 16'h9c2b, 16'h99f1, 16'h99cb,
// 16'h9bb2, 16'h9fa9, 16'ha58b, 16'had4b,
// 16'hb6b1, 16'hc198, 16'hcdbf, 16'hdaef,
// 16'he8da, 16'hf744, 16'h05d4, 16'h144a,
// 16'h2257, 16'h2fae, 16'h3c15, 16'h473b,
// 16'h50f7, 16'h590a, 16'h5f53, 16'h63ab,
// 16'h65fe, 16'h6642, 16'h6470, 16'h6098,
// 16'h5aca, 16'h5324, 16'h49d1, 16'h3efb,
// 16'h32e4, 16'h25be, 16'h17dc, 16'h0977,
// 16'hfae6, 16'hec6d, 16'hde59, 16'hd0f7,
// 16'hc484, 16'hb94b, 16'haf7c, 16'ha752,
// 16'ha0f2, 16'h9c82, 16'h9a11, 16'h99b7,
// 16'h9b6b, 16'h9f2b, 16'ha4e0, 16'hac70,
// 16'hb5ad, 16'hc074, 16'hcc79, 16'hd995,
// 16'he76f, 16'hf5ce, 16'h0462, 16'h12d8,
// 16'h20f9, 16'h2e62, 16'h3ae3, 16'h4630,
// 16'h500c, 16'h5854, 16'h5ec5, 16'h6353,
// 16'h65dd, 16'h664e, 16'h64bb, 16'h6110,
// 16'h5b73, 16'h53ff, 16'h4acd, 16'h4025,
// 16'h3423, 16'h271b, 16'h1944, 16'h0aec,
// 16'hfc5b, 16'heddc, 16'hdfbb, 16'hd243,
// 16'hc5b6, 16'hba5c, 16'hb063, 16'ha811,
// 16'ha17f, 16'h9cdb, 16'h9a3b, 16'h99a4,
// 16'h9b2b, 16'h9eb1, 16'ha43c, 16'hab96,
// 16'hb4b2, 16'hbf4c, 16'hcb3c, 16'hd839,
// 16'he606, 16'hf45c, 16'h02e9, 16'h116e,
// 16'h1f92, 16'h2d16, 16'h39b0, 16'h451c,
// 16'h4f25, 16'h5790, 16'h5e39, 16'h62f4,
// 16'h65b2, 16'h665f, 16'h64f5, 16'h618a,
// 16'h5c15, 16'h54d5, 16'h4bc9, 16'h4146,
// 16'h3564, 16'h2872, 16'h1aaf, 16'h0c5e,
// 16'hfdd0, 16'hef4d, 16'he11e, 16'hd392,
// 16'hc6ec, 16'hbb6d, 16'hb154, 16'ha8ce,
// 16'ha215, 16'h9d38, 16'h9a69, 16'h999a,
// 16'h9aed, 16'h9e3f, 16'ha398, 16'haac6,
// 16'hb3b7, 16'hbe2b, 16'hc9fe, 16'hd6e1,
// 16'he49f, 16'hf2e8, 16'h0175, 16'h0ffc,
// 16'h1e2d, 16'h2bc9, 16'h3875, 16'h440c,
// 16'h4e32, 16'h56ce, 16'h5da4, 16'h6291,
// 16'h6584, 16'h6665, 16'h6533, 16'h61f5,
// 16'h5cbb, 16'h559e, 16'h4cc8, 16'h4262,
// 16'h36a0, 16'h29ca, 16'h1c15, 16'h0dd2,
// 16'hff45, 16'hf0bd, 16'he284, 16'hd4e3,
// 16'hc825, 16'hbc82, 16'hb245, 16'ha996,
// 16'ha2aa, 16'h9da0, 16'h9a98, 16'h9997,
// 16'h9ab2, 16'h9dd5, 16'ha2f6, 16'ha9fe,
// 16'hb2ba, 16'hbd15, 16'hc8bd, 16'hd58f,
// 16'he337, 16'hf174, 16'h2002, 16'h0e89,
// 16'h1cca, 16'h2a72, 16'h3740, 16'h42ef,
// 16'h4d42, 16'h5606, 16'h5d06, 16'h622e,
// 16'h654d, 16'h6668, 16'h6569, 16'h6261,
// 16'h5d53, 16'h566e, 16'h4db8, 16'h437e,
// 16'h37dd, 16'h2b1b, 16'h1d7e, 16'h0f41,
// 16'h20bd, 16'hf22c, 16'he3ed, 16'hd635,
// 16'hc960, 16'hbd9d, 16'hb33b, 16'haa5f,
// 16'ha347, 16'h9e0a, 16'h9acd, 16'h999b,
// 16'h9a7c, 16'h9d6f, 16'ha25c, 16'ha934,
// 16'hb1ca, 16'hbbf8, 16'hc787, 16'hd43c,
// 16'he1cf, 16'hf007, 16'hfe88, 16'h0d1a,
// 16'h1b60, 16'h2920, 16'h3602, 16'h41d4,
// 16'h4c4a, 16'h5538, 16'h5c6c, 16'h61bc,
// 16'h6517, 16'h6663, 16'h659a, 16'h62c6,
// 16'h5ded, 16'h572f, 16'h4eae, 16'h4492,
// 16'h3915, 16'h2c6e, 16'h1ee1, 16'h10b5,
// 16'h022d, 16'hf3a5, 16'he54f, 16'hd790,
// 16'hca9a, 16'hbebc, 16'hb434, 16'hab2e,
// 16'ha3e9, 16'h9e78, 16'h9b09, 16'h99a2,
// 16'h9a4d, 16'h9d0d, 16'ha1c7, 16'ha870,
// 16'hb0da, 16'hbae4, 16'hc651, 16'hd2ea,
// 16'he06e, 16'hee92, 16'hfd16, 16'h0ba6,
// 16'h19f7, 16'h27cb, 16'h34c1, 16'h40b6,
// 16'h4b4d, 16'h5468, 16'h5bc7, 16'h614d,
// 16'h64d8, 16'h6658, 16'h65c8, 16'h6324,
// 16'h5e7f, 16'h57f4, 16'h4f98, 16'h45a7,
// 16'h3a4b, 16'h2db9, 16'h2049, 16'h1220,
// 16'h03a9, 16'hf511, 16'he6be, 16'hd8e3,
// 16'hcbde, 16'hbfdc, 16'hb531, 16'hac02,
// 16'ha48d, 16'h9eef, 16'h9b48, 16'h99af,
// 16'h9a23, 16'h9cb0, 16'ha137, 16'ha7b0,
// 16'haff1, 16'hb9d1, 16'hc51e, 16'hd19c,
// 16'hdf0a, 16'hed24, 16'hfba1, 16'h0a32,
// 16'h1890, 16'h266c, 16'h3384, 16'h3f91,
// 16'h4a4f, 16'h5393, 16'h5b1e, 16'h60d5,
// 16'h6497, 16'h6646, 16'h65f3, 16'h637a,
// 16'h5f12, 16'h58ab, 16'h5085, 16'h46b5,
// 16'h3b7c, 16'h2f0a, 16'h21a4, 16'h1397,
// 16'h0516, 16'hf68c, 16'he824, 16'hda3f,
// 16'hcd20, 16'hc101, 16'hb633, 16'hacda,
// 16'ha536, 16'h9f69, 16'h9b8e, 16'h99c0,
// 16'h9a02, 16'h9c53, 16'ha0b0, 16'ha6f3,
// 16'haf0b, 16'hb8c3, 16'hc3ee, 16'hd04f,
// 16'hddab, 16'hebb5, 16'hfa2b, 16'h08be,
// 16'h1725, 16'h2510, 16'h3244, 16'h3e63,
// 16'h4954, 16'h52b2, 16'h5a77, 16'h6056,
// 16'h644e, 16'h6634, 16'h6612, 16'h63d2,
// 16'h5f98, 16'h5966, 16'h5167, 16'h47c4,
// 16'h3ca9, 16'h3053, 16'h2309, 16'h14fe,
// 16'h0691, 16'hf7fc, 16'he991, 16'hdb9d,
// 16'hce63, 16'hc22b, 16'hb735, 16'hadb7,
// 16'ha5e7, 16'h9fe5, 16'h9bdd, 16'h99d2,
// 16'h99e6, 16'h9c20, 16'ha029, 16'ha63e,
// 16'hae28, 16'hb7b8, 16'hc2c2, 16'hcf05,
// 16'hdc4d, 16'hea47, 16'hf8b6, 16'h074b,
// 16'h15b6, 16'h23b7, 16'h30f8, 16'h3d3f,
// 16'h4848, 16'h51d8, 16'h59c2, 16'h5fd8,
// 16'h63fd, 16'h661e, 16'h662a, 16'h6425,
// 16'h601b, 16'h5a19, 16'h5249, 16'h48cb,
// 16'h3dd4, 16'h319d, 16'h2464, 16'h166e,
// 16'h0804, 16'hf971, 16'heafe, 16'hdcfb,
// 16'hcfaa, 16'hc358, 16'hb83d, 16'hae98,
// 16'ha69a, 16'ha06a, 16'h9c29, 16'h99f5,
// 16'h99c6, 16'h9bb7, 16'h9fa6, 16'ha58c,
// 16'had4b, 16'hb6b0, 16'hc199, 16'hcdbf,
// 16'hdaee, 16'he8dc, 16'hf741, 16'h05d6,
// 16'h144b, 16'h2254, 16'h2fb2, 16'h3c10,
// 16'h473f, 16'h50f5, 16'h590c, 16'h5f51,
// 16'h63ac, 16'h65fe, 16'h6641, 16'h6472,
// 16'h6096, 16'h5acb, 16'h5325, 16'h49ce,
// 16'h3eff, 16'h32e0, 16'h25c1, 16'h17da,
// 16'h0978, 16'hfae6, 16'hec6c, 16'hde5b,
// 16'hd0f4, 16'hc487, 16'hb949, 16'haf7d,
// 16'ha752, 16'ha0f2, 16'h9c81, 16'h9a12,
// 16'h99b7, 16'h9b6a, 16'h9f2d, 16'ha4de,
// 16'hac71, 16'hb5ae, 16'hc072, 16'hcc7a,
// 16'hd995, 16'he76e, 16'hf5d1, 16'h045d,
// 16'h12dd, 16'h20f5, 16'h2e64, 16'h3ae4,
// 16'h462c, 16'h5011, 16'h5850, 16'h5ec7,
// 16'h6354, 16'h65d9, 16'h6654, 16'h64b6,
// 16'h6112, 16'h5b73, 16'h53fe, 16'h4ad0,
// 16'h4021, 16'h3427, 16'h2717, 16'h1947,
// 16'h0aeb, 16'hfc5a, 16'hedde, 16'hdfb9,
// 16'hd245, 16'hc5b4, 16'hba5d, 16'hb063,
// 16'ha810, 16'ha181, 16'h9cd9, 16'h9a3b,
// 16'h99a7, 16'h9b26, 16'h9eb7, 16'ha436,
// 16'hab9a, 16'hb4b0, 16'hbf4d, 16'hcb3c,
// 16'hd837, 16'he609, 16'hf459, 16'h02eb,
// 16'h116d, 16'h1f91, 16'h2d18, 16'h39ae,
// 16'h451d, 16'h4f26, 16'h578e, 16'h5e3a,
// 16'h62f3, 16'h65b4, 16'h665c, 16'h64fa,
// 16'h6184, 16'h5c1b, 16'h54cf, 16'h4bcf,
// 16'h4141, 16'h3568, 16'h286f, 16'h1ab1,
// 16'h0c5d, 16'hfdd0, 16'hef4c, 16'he120,
// 16'hd38f, 16'hc6f0, 16'hbb68, 16'hb157,
// 16'ha8cf, 16'ha211, 16'h9d3e, 16'h9a62,
// 16'h99a0, 16'h9ae9, 16'h9e42, 16'ha395,
// 16'haac9, 16'hb3b3, 16'hbe30, 16'hc9fa,
// 16'hd6e4, 16'he49c, 16'hf2ea, 16'h0174,
// 16'h0ffc, 16'h1e2f, 16'h2bc5, 16'h387a,
// 16'h4408, 16'h4e34, 16'h56cd, 16'h5da4,
// 16'h6291, 16'h6586, 16'h6661, 16'h6538,
// 16'h61f0, 16'h5cbf, 16'h559c, 16'h4cc9,
// 16'h4260, 16'h36a3, 16'h29c7, 16'h1c17,
// 16'h0dd1, 16'hff46, 16'hf0bc, 16'he285,
// 16'hd4e2, 16'hc824, 16'hbc85, 16'hb243,
// 16'ha997, 16'ha2a9, 16'h9da1, 16'h9a96,
// 16'h999a, 16'h9ab0, 16'h9dd6, 16'ha2f6,
// 16'ha9fc, 16'hb2be, 16'hbd10, 16'hc8c2,
// 16'hd58b, 16'he339, 16'hf174, 16'h2001,
// 16'h0e8a, 16'h1cc9, 16'h2a73, 16'h373f,
// 16'h42f0, 16'h4d41, 16'h5606, 16'h5d08,
// 16'h622c, 16'h654e, 16'h6668, 16'h6568,
// 16'h6261, 16'h5d55, 16'h566b, 16'h4dbb,
// 16'h437d, 16'h37da, 16'h2b20, 16'h1d78,
// 16'h0f47, 16'h20b8, 16'hf230, 16'he3ea,
// 16'hd637, 16'hc95d, 16'hbda1, 16'hb337,
// 16'haa63, 16'ha344, 16'h9e0b, 16'h9acd,
// 16'h999c, 16'h9a7a, 16'h9d72, 16'ha258,
// 16'ha937, 16'hb1c9, 16'hbbf8, 16'hc788,
// 16'hd43b, 16'he1cf, 16'hf007, 16'hfe89,
// 16'h0d19, 16'h1b62, 16'h291d, 16'h3605,
// 16'h41d2, 16'h4c4b, 16'h5539, 16'h5c68,
// 16'h61c1, 16'h6514, 16'h6664, 16'h659a,
// 16'h62c5, 16'h5ded, 16'h5731, 16'h4eac,
// 16'h4493, 16'h3915, 16'h2c6d, 16'h1ee2,
// 16'h10b4, 16'h022f, 16'hf3a2, 16'he551,
// 16'hd790, 16'hca98, 16'hbec0, 16'hb42f,
// 16'hab33, 16'ha3e4, 16'h9e7d, 16'h9b05,
// 16'h99a4, 16'h9a4d, 16'h9d0b, 16'ha1c9,
// 16'ha86e, 16'hb0dd, 16'hbae2, 16'hc651,
// 16'hd2ea, 16'he06d, 16'hee94, 16'hfd16,
// 16'h0ba4, 16'h19fb, 16'h27c5, 16'h34c7,
// 16'h40b1, 16'h4b51, 16'h5466, 16'h5bc8,
// 16'h614c, 16'h64d7, 16'h665b, 16'h65c5,
// 16'h6325, 16'h5e81, 16'h57f0, 16'h4f9b,
// 16'h45a7, 16'h3a47, 16'h2dbf, 16'h2044,
// 16'h1224, 16'h03a6, 16'hf513, 16'he6bc,
// 16'hd8e5, 16'hcbdc, 16'hbfde, 16'hb530,
// 16'hac02, 16'ha48e, 16'h9eed, 16'h9b4a,
// 16'h99ad, 16'h9a25, 16'h9caf, 16'ha137,
// 16'ha7b0, 16'haff2, 16'hb9cf, 16'hc520,
// 16'hd19a, 16'hdf0c, 16'hed24, 16'hfba0,
// 16'h0a32, 16'h188f, 16'h266e, 16'h3384,
// 16'h3f8f, 16'h4a52, 16'h538f, 16'h5b22,
// 16'h60d2, 16'h6498, 16'h6648, 16'h65ee,
// 16'h6381, 16'h5f0a, 16'h58b2, 16'h5080,
// 16'h46b9, 16'h3b79, 16'h2f0a, 16'h21a7,
// 16'h1393, 16'h051a, 16'hf689, 16'he824,
// 16'hda42, 16'hcd1d, 16'hc104, 16'hb630,
// 16'hacda, 16'ha539, 16'h9f65, 16'h9b93,
// 16'h99bb, 16'h9a04, 16'h9c53, 16'ha0b0,
// 16'ha6f3, 16'haf0a, 16'hb8c5, 16'hc3eb,
// 16'hd053, 16'hdda7, 16'hebb8, 16'hfa2a,
// 16'h08bf, 16'h1723, 16'h2513, 16'h323f,
// 16'h3e6b, 16'h494b, 16'h52ba, 16'h5a70,
// 16'h605b, 16'h644b, 16'h6637, 16'h660e,
// 16'h63d5, 16'h5f96, 16'h5967, 16'h5168,
// 16'h47c1, 16'h3cab, 16'h3052, 16'h2309,
// 16'h1520, 16'h068f, 16'hf7fd, 16'he990,
// 16'hdb9e, 16'hce62, 16'hc22d, 16'hb734,
// 16'hadb8, 16'ha5e6, 16'h9fe5, 16'h9bdd,
// 16'h99d3, 16'h99e5, 16'h9c20, 16'ha02a,
// 16'ha63d, 16'hae28, 16'hb7b9, 16'hc2bf,
// 16'hcf09, 16'hdc4a, 16'hea48, 16'hf8b7,
// 16'h0749, 16'h15b8, 16'h23b5, 16'h30f9,
// 16'h3d40, 16'h4846, 16'h51db, 16'h59bd,
// 16'h5fde, 16'h63f8, 16'h6622, 16'h6627,
// 16'h6428, 16'h6018, 16'h5a1c, 16'h5246,
// 16'h48ce, 16'h3dd1, 16'h31a0, 16'h2461,
// 16'h1671, 16'h0802, 16'hf971, 16'heaff,
// 16'hdcfa, 16'hcfab, 16'hc358, 16'hb83c,
// 16'hae98, 16'ha69b, 16'ha068, 16'h9c2d,
// 16'h99f0, 16'h99ca, 16'h9bb3, 16'h9faa,
// 16'ha589, 16'had4d, 16'hb6af, 16'hc199,
// 16'hcdc0, 16'hdaec, 16'he8df, 16'hf73d,
// 16'h05da, 16'h1447, 16'h2258, 16'h2faf,
// 16'h3c12, 16'h473c, 16'h50f9, 16'h5908,
// 16'h5f55, 16'h63a8, 16'h6620, 16'h6642,
// 16'h646f, 16'h609a, 16'h5ac7, 16'h5327,
// 16'h49ce, 16'h3efe, 16'h32e1, 16'h25c1,
// 16'h17d9, 16'h097a, 16'hfae3, 16'hec6f,
// 16'hde58, 16'hd0f7, 16'hc485, 16'hb94a,
// 16'haf7d, 16'ha751, 16'ha0f3, 16'h9c80,
// 16'h9a14, 16'h99b4, 16'h9b6d, 16'h9f2a,
// 16'ha4e0, 16'hac70, 16'hb5ae, 16'hc072,
// 16'hcc7b, 16'hd993, 16'he770, 16'hf5cf,
// 16'h045f, 16'h12dc, 16'h20f6, 16'h2e63,
// 16'h3ae4, 16'h462d, 16'h5010, 16'h5851,
// 16'h5ec6, 16'h6355, 16'h65d7, 16'h6656,
// 16'h64b4, 16'h6114, 16'h5b73, 16'h53fb,
// 16'h4ad3, 16'h4020, 16'h3425, 16'h271b,
// 16'h1944, 16'h0aec, 16'hfc5b, 16'heddb,
// 16'hdfbc, 16'hd243, 16'hc5b7, 16'hba59,
// 16'hb067, 16'ha80c, 16'ha183, 16'h9cd9,
// 16'h9a3b, 16'h99a6, 16'h9b28, 16'h9eb4,
// 16'ha439, 16'hab98, 16'hb4b2, 16'hbf4b,
// 16'hcb3d, 16'hd838, 16'he608, 16'hf459,
// 16'h02ec, 16'h116b, 16'h1f93, 16'h2d17,
// 16'h39ae, 16'h451e, 16'h4f24, 16'h578f,
// 16'h5e3b, 16'h62f2, 16'h65b4, 16'h665d,
// 16'h64f7, 16'h6188, 16'h5c17, 16'h54d2,
// 16'h4bcd, 16'h4143, 16'h3566, 16'h2870,
// 16'h1ab1, 16'h0c5d, 16'hfdd0, 16'hef4d,
// 16'he11e, 16'hd392, 16'hc6ec, 16'hbb6d,
// 16'hb152, 16'ha8d3, 16'ha20f, 16'h9d3d,
// 16'h9a64, 16'h999f, 16'h9ae9, 16'h9e42,
// 16'ha395, 16'haac9, 16'hb3b3, 16'hbe31,
// 16'hc9f8, 16'hd6e6, 16'he49c, 16'hf2e8,
// 16'h0175, 16'h0ffd, 16'h1e2e, 16'h2bc5,
// 16'h387b, 16'h4404, 16'h4e39, 16'h56cb,
// 16'h5da3, 16'h6293, 16'h6583, 16'h6665,
// 16'h6533, 16'h61f6, 16'h5cb9, 16'h55a1,
// 16'h4cc4, 16'h4265, 16'h369e, 16'h29cc,
// 16'h1c14, 16'h0dd1, 16'hff48, 16'hf0b9,
// 16'he287, 16'hd4e2, 16'hc825, 16'hbc83,
// 16'hb244, 16'ha996, 16'ha2ab, 16'h9d9f,
// 16'h9a97, 16'h999a, 16'h9aaf, 16'h9dd8,
// 16'ha2f4, 16'ha9fd, 16'hb2bc, 16'hbd14,
// 16'hc8bd, 16'hd591, 16'he334, 16'hf176,
// 16'h2002, 16'h0e87, 16'h1ccc, 16'h2a72,
// 16'h373f, 16'h42f1, 16'h4d3f, 16'h5608,
// 16'h5d05, 16'h6230, 16'h654b, 16'h6669,
// 16'h6569, 16'h625f, 16'h5d57, 16'h566a,
// 16'h4dbb, 16'h437c, 16'h37dd, 16'h2b1d,
// 16'h1d7b, 16'h0f45, 16'h20b7, 16'hf232,
// 16'he3e9, 16'hd638, 16'hc95e, 16'hbd9d,
// 16'hb33c, 16'haa5e, 16'ha349, 16'h9e08,
// 16'h9acd, 16'h999d, 16'h9a7a, 16'h9d70,
// 16'ha25c, 16'ha932, 16'hb1cd, 16'hbbf6,
// 16'hc789, 16'hd43a, 16'he1cf, 16'hf008,
// 16'hfe87, 16'h0d1c, 16'h1b5f, 16'h291f,
// 16'h3604, 16'h41d1, 16'h4c4d, 16'h5536,
// 16'h5c6c, 16'h61be, 16'h6515, 16'h6663,
// 16'h659b, 16'h62c4, 16'h5def, 16'h572e,
// 16'h4eae, 16'h4493, 16'h3913, 16'h2c70,
// 16'h1ee0, 16'h10b4, 16'h0230, 16'hf3a2,
// 16'he551, 16'hd78f, 16'hca99, 16'hbebf,
// 16'hb431, 16'hab31, 16'ha3e5, 16'h9e7c,
// 16'h9b06, 16'h99a4, 16'h9a4d, 16'h9d0b,
// 16'ha1c8, 16'ha870, 16'hb0db, 16'hbae3,
// 16'hc652, 16'hd2e8, 16'he06f, 16'hee93,
// 16'hfd15, 16'h0ba6, 16'h19f9, 16'h27c7,
// 16'h34c6, 16'h40b1, 16'h4b51, 16'h5466,
// 16'h5bc7, 16'h614e, 16'h64d7, 16'h6658,
// 16'h65c9, 16'h6321, 16'h5e84, 16'h57ee,
// 16'h4f9d, 16'h45a4, 16'h3a4b, 16'h2dbc,
// 16'h2044, 16'h1226, 16'h03a3, 16'hf516,
// 16'he6bb, 16'hd8e5, 16'hcbdc, 16'hbfde,
// 16'hb52f, 16'hac04, 16'ha48c, 16'h9eee,
// 16'h9b4a, 16'h99ac, 16'h9a28, 16'h9caa,
// 16'ha13b, 16'ha7ae, 16'haff2, 16'hb9d1,
// 16'hc51d, 16'hd19c, 16'hdf0b, 16'hed24,
// 16'hfba1, 16'h0a30, 16'h1891, 16'h266d,
// 16'h3384, 16'h3f90, 16'h4a50, 16'h5391,
// 16'h5b20, 16'h60d4, 16'h6497, 16'h6648,
// 16'h65ef, 16'h637d, 16'h5f10, 16'h58ad,
// 16'h5083, 16'h46b8, 16'h3b78, 16'h2f0c,
// 16'h21a5, 16'h1394, 16'h051a, 16'hf689,
// 16'he824, 16'hda42, 16'hcd1b, 16'hc106,
// 16'hb62f, 16'hacdb, 16'ha538, 16'h9f66,
// 16'h9b91, 16'h99be, 16'h9a01, 16'h9c55,
// 16'ha0b0, 16'ha6f1, 16'haf0f, 16'hb8be,
// 16'hc3f1, 16'hd04f, 16'hddab, 16'hebb4,
// 16'hfa2d, 16'h08bc, 16'h1726, 16'h2512,
// 16'h323f, 16'h3e6b, 16'h494a, 16'h52bd,
// 16'h5a6c, 16'h605f, 16'h6449, 16'h6636,
// 16'h6610, 16'h63d4, 16'h5f97, 16'h5966,
// 16'h5168, 16'h47c1, 16'h3cac, 16'h3052,
// 16'h2309, 16'h14fe, 16'h0692, 16'hf7fa,
// 16'he993, 16'hdb9c, 16'hce63, 16'hc22c,
// 16'hb734, 16'hadb8, 16'ha5e7, 16'h9fe3,
// 16'h9bdf, 16'h99d1, 16'h99e7, 16'h9bff,
// 16'ha02a, 16'ha63d, 16'hae28, 16'hb7ba,
// 16'hc2be, 16'hcf0a, 16'hdc49, 16'hea48,
// 16'hf8b8, 16'h0748, 16'h15b9, 16'h23b4,
// 16'h30fa, 16'h3d3f, 16'h4848, 16'h51d7,
// 16'h59c3, 16'h5fd6, 16'h6401, 16'h661b,
// 16'h662b, 16'h6426, 16'h6018, 16'h5a1c,
// 16'h5248, 16'h48ca, 16'h3dd7, 16'h3199,
// 16'h2468, 16'h166b, 16'h0806, 16'hf96f,
// 16'heb20, 16'hdcfa, 16'hcfab, 16'hc357,
// 16'hb83d, 16'hae98, 16'ha69a, 16'ha06a,
// 16'h9c2a, 16'h99f3, 16'h99c8, 16'h9bb5,
// 16'h9fa6, 16'ha58e, 16'had49, 16'hb6b2,
// 16'hc197, 16'hcdc0, 16'hdaed, 16'he8de,
// 16'hf740, 16'h05d5, 16'h144c, 16'h2253,
// 16'h2fb4, 16'h3c0e, 16'h4741, 16'h50f3,
// 16'h590c, 16'h5f53, 16'h63a9, 16'h6601,
// 16'h6640, 16'h6470, 16'h609a, 16'h5ac6,
// 16'h5329, 16'h49cb, 16'h3f02, 16'h32de,
// 16'h25c3, 16'h17d7, 16'h097b, 16'hfae4,
// 16'hec6d, 16'hde5b, 16'hd0f4, 16'hc487,
// 16'hb949, 16'haf7d, 16'ha752, 16'ha0f2,
// 16'h9c81, 16'h9a12, 16'h99b7, 16'h9b6b,
// 16'h9f2a, 16'ha4e2, 16'hac6d, 16'hb5b1,
// 16'hc06f, 16'hcc7d, 16'hd993, 16'he76f,
// 16'hf5d0, 16'h045e, 16'h12dd, 16'h20f4,
// 16'h2e66, 16'h3ae1, 16'h4630, 16'h500e,
// 16'h5851, 16'h5ec7, 16'h6353, 16'h65da,
// 16'h6653, 16'h64b7, 16'h6111, 16'h5b74,
// 16'h53fc, 16'h4ad1, 16'h4022, 16'h3424,
// 16'h271c, 16'h1942, 16'h0aef, 16'hfc57,
// 16'heddf, 16'hdfba, 16'hd244, 16'hc5b6,
// 16'hba5a, 16'hb065, 16'ha80f, 16'ha180,
// 16'h9cdc, 16'h9a38, 16'h99a9, 16'h9b25,
// 16'h9eb7, 16'ha436, 16'hab9b, 16'hb4b0,
// 16'hbf4c, 16'hcb3d, 16'hd837, 16'he609,
// 16'hf458, 16'h02ed, 16'h116a, 16'h1f95,
// 16'h2d14, 16'h39b1, 16'h451b, 16'h4f25,
// 16'h5792, 16'h5e36, 16'h62f7, 16'h65af,
// 16'h6661, 16'h64f5, 16'h6189, 16'h5c16,
// 16'h54d4, 16'h4bca, 16'h4146, 16'h3563,
// 16'h2873, 16'h1aaf, 16'h0c5d, 16'hfdd1,
// 16'hef4c, 16'he11e, 16'hd394, 16'hc6ea,
// 16'hbb6d, 16'hb154, 16'ha8ce, 16'ha216,
// 16'h9d38, 16'h9a67, 16'h999d, 16'h9ae9,
// 16'h9e44, 16'ha394, 16'haac8, 16'hb3b5,
// 16'hbe2e, 16'hc9fb, 16'hd6e5, 16'he49b,
// 16'hf2ea, 16'h0173, 16'h0ffd, 16'h1e2f,
// 16'h2bc5, 16'h387a, 16'h4406, 16'h4e36,
// 16'h56cd, 16'h5da4, 16'h6291, 16'h6585,
// 16'h6662, 16'h6536, 16'h61f5, 16'h5cba,
// 16'h559f, 16'h4cc7, 16'h4260, 16'h36a4,
// 16'h29c8, 16'h1c16, 16'h0dd0, 16'hff47,
// 16'hf0bb, 16'he287, 16'hd4e0, 16'hc826,
// 16'hbc82, 16'hb246, 16'ha995, 16'ha2aa,
// 16'h9da1, 16'h9a95, 16'h999b, 16'h9ab0,
// 16'h9dd5, 16'ha2f7, 16'ha9fc, 16'hb2bc,
// 16'hbd14, 16'hc8bd, 16'hd590, 16'he335,
// 16'hf177, 16'hffff, 16'h0e8b, 16'h1cc8,
// 16'h2a75, 16'h373d, 16'h42f1, 16'h4d41,
// 16'h5605, 16'h5d0a, 16'h622a, 16'h654f,
// 16'h6668, 16'h6567, 16'h6263, 16'h5d54,
// 16'h566a, 16'h4dbd, 16'h437a, 16'h37df,
// 16'h2b1a, 16'h1d7f, 16'h0f3f, 16'h20bf,
// 16'hf22b, 16'he3ed, 16'hd636, 16'hc95e,
// 16'hbd9f, 16'hb339, 16'haa61, 16'ha345,
// 16'h9e0c, 16'h9acb, 16'h999d, 16'h9a7b,
// 16'h9d6f, 16'ha25c, 16'ha934, 16'hb1ca,
// 16'hbbf8, 16'hc789, 16'hd438, 16'he1d3,
// 16'hf004, 16'hfe89, 16'h0d1a, 16'h1b62,
// 16'h291b, 16'h3608, 16'h41cf, 16'h4c4d,
// 16'h5538, 16'h5c68, 16'h61c2, 16'h6513,
// 16'h6665, 16'h6599, 16'h62c6, 16'h5dec,
// 16'h5731, 16'h4ead, 16'h4493, 16'h3915,
// 16'h2c6d, 16'h1ee1, 16'h10b4, 16'h0232,
// 16'hf39e, 16'he555, 16'hd78c, 16'hca9b,
// 16'hbebe, 16'hb431, 16'hab30, 16'ha3e9,
// 16'h9e76, 16'h9b0c, 16'h999f, 16'h9a50,
// 16'h9d0a, 16'ha1c9, 16'ha86e, 16'hb0dd,
// 16'hbae2, 16'hc652, 16'hd2e9, 16'he06e,
// 16'hee93, 16'hfd16, 16'h0ba6, 16'h19f8,
// 16'h27c8, 16'h34c5, 16'h40b2, 16'h4b51,
// 16'h5465, 16'h5bc9, 16'h614b, 16'h64da,
// 16'h6656, 16'h65ca, 16'h6321, 16'h5e83,
// 16'h57f0, 16'h4f9a, 16'h45a7, 16'h3a48,
// 16'h2dbe, 16'h2045, 16'h1222, 16'h03a7,
// 16'hf513, 16'he6be, 16'hd8e3, 16'hcbdd,
// 16'hbfdc, 16'hb532, 16'hac02, 16'ha48d,
// 16'h9eee, 16'h9b49, 16'h99ae, 16'h9a25,
// 16'h9cad, 16'ha13a, 16'ha7ae, 16'haff2,
// 16'hb9d0, 16'hc51f, 16'hd19b, 16'hdf0b,
// 16'hed25, 16'hfb9e, 16'h0a35, 16'h188c,
// 16'h2671, 16'h3381, 16'h3f91, 16'h4a50,
// 16'h5392, 16'h5b1e, 16'h60d7, 16'h6493,
// 16'h664b, 16'h65ee, 16'h637d, 16'h5f11,
// 16'h58ab, 16'h5086, 16'h46b4, 16'h3b7c,
// 16'h2f0a, 16'h21a5, 16'h1394, 16'h051b,
// 16'hf686, 16'he829, 16'hda3c, 16'hcd21,
// 16'hc102, 16'hb630, 16'hacdc, 16'ha535,
// 16'h9f6b, 16'h9b8b, 16'h99c4, 16'h99fc,
// 16'h9c59, 16'ha0ab, 16'ha6f7, 16'haf09,
// 16'hb8c4, 16'hc3ec, 16'hd052, 16'hdda8,
// 16'hebb8, 16'hfa29, 16'h08bf, 16'h1725,
// 16'h2510, 16'h3242, 16'h3e67, 16'h4950,
// 16'h52b5, 16'h5a75, 16'h6057, 16'h644d,
// 16'h6636, 16'h660f, 16'h63d5, 16'h5f96,
// 16'h5967, 16'h5167, 16'h47c4, 16'h3ca7,
// 16'h3057, 16'h2305, 16'h1501, 16'h0691,
// 16'hf7fa, 16'he992, 16'hdb9f, 16'hce5e,
// 16'hc231, 16'hb732, 16'hadb7, 16'ha5e9,
// 16'h9fe2, 16'h9bde, 16'h99d4, 16'h99e3,
// 16'h9c03, 16'ha026, 16'ha641, 16'hae25,
// 16'hb7bb, 16'hc2bf, 16'hcf08, 16'hdc4b,
// 16'hea46, 16'hf8b9, 16'h0747, 16'h15bb,
// 16'h23b2, 16'h30fb, 16'h3d3d, 16'h484a,
// 16'h51d6, 16'h59c4, 16'h5fd5, 16'h6402,
// 16'h6618, 16'h6630, 16'h6421, 16'h601d,
// 16'h5a18, 16'h5249, 16'h48cc, 16'h3dd3,
// 16'h319e, 16'h2463, 16'h166e, 16'h0805,
// 16'hf970, 16'heaff, 16'hdcfa, 16'hcfab,
// 16'hc357, 16'hb83e, 16'hae98, 16'ha699,
// 16'ha06a, 16'h9c2b, 16'h99f1, 16'h99cb,
// 16'h9bb3, 16'h9fa7, 16'ha58d, 16'had49,
// 16'hb6b3, 16'hc196, 16'hcdc1, 16'hdaed,
// 16'he8dc, 16'hf742, 16'h05d6, 16'h1448,
// 16'h2259, 16'h2fad, 16'h3c15, 16'h473b,
// 16'h50f7, 16'h590b, 16'h5f52, 16'h63ac,
// 16'h65fd, 16'h6642, 16'h6471, 16'h6098,
// 16'h5aca, 16'h5323, 16'h49d2, 16'h3efa,
// 16'h32e6, 16'h25bc, 16'h17dd, 16'h0976,
// 16'hfae7, 16'hec6c, 16'hde5b, 16'hd0f4,
// 16'hc486, 16'hb94b, 16'haf7a, 16'ha756,
// 16'ha0ee, 16'h9c84, 16'h9a10, 16'h99b9,
// 16'h9b67, 16'h9f30, 16'ha4db, 16'hac74,
// 16'hb5ac, 16'hc071, 16'hcc7e, 16'hd990,
// 16'he773, 16'hf5cc, 16'h0461, 16'h12dc,
// 16'h20f4, 16'h2e67, 16'h3ade, 16'h4634,
// 16'h500b, 16'h5853, 16'h5ec5, 16'h6355,
// 16'h65d9, 16'h6654, 16'h64b6, 16'h6111,
// 16'h5b75, 16'h53fc, 16'h4ad1, 16'h4021,
// 16'h3426, 16'h2719, 16'h1946, 16'h0aea,
// 16'hfc5d, 16'hedd9, 16'hdfbf, 16'hd23f,
// 16'hc5bb, 16'hba56, 16'hb069, 16'ha80b,
// 16'ha184, 16'h9cd8, 16'h9a3b, 16'h99a7,
// 16'h9b27, 16'h9eb5, 16'ha437, 16'hab9a,
// 16'hb4b1, 16'hbf4b, 16'hcb3e, 16'hd836,
// 16'he609, 16'hf45a, 16'h02eb, 16'h116b,
// 16'h1f94, 16'h2d16, 16'h39ae, 16'h451f,
// 16'h4f22, 16'h5793, 16'h5e36, 16'h62f7,
// 16'h65b0, 16'h665f, 16'h64f8, 16'h6185,
// 16'h5c1b, 16'h54cf, 16'h4bce, 16'h4143,
// 16'h3565, 16'h2872, 16'h1aaf, 16'h0c5e,
// 16'hfdd0, 16'hef4d, 16'he11d, 16'hd393,
// 16'hc6ed, 16'hbb6a, 16'hb157, 16'ha8cc,
// 16'ha215, 16'h9d3b, 16'h9a64, 16'h999f,
// 16'h9ae9, 16'h9e41, 16'ha398, 16'haac5,
// 16'hb3b8, 16'hbe2b, 16'hc9fe, 16'hd6e1,
// 16'he49e, 16'hf2e9, 16'h0173, 16'h1020,
// 16'h1e29, 16'h2bcb, 16'h3874, 16'h440c,
// 16'h4e31, 16'h56d1, 16'h5da0, 16'h6294,
// 16'h6583, 16'h6664, 16'h6535, 16'h61f3,
// 16'h5cbd, 16'h559d, 16'h4cc9, 16'h425f,
// 16'h36a3, 16'h29c9, 16'h1c15, 16'h0dd3,
// 16'hff43, 16'hf0bf, 16'he281, 16'hd4e6,
// 16'hc822, 16'hbc85, 16'hb244, 16'ha996,
// 16'ha2a8, 16'h9da3, 16'h9a94, 16'h999c,
// 16'h9ab0, 16'h9dd4, 16'ha2f8, 16'ha9fa,
// 16'hb2bf, 16'hbd11, 16'hc8c0, 16'hd58d,
// 16'he337, 16'hf176, 16'hffff, 16'h0e8c,
// 16'h1cc7, 16'h2a75, 16'h373e, 16'h42f0,
// 16'h4d42, 16'h5604, 16'h5d0b, 16'h6228,
// 16'h6552, 16'h6665, 16'h656a, 16'h6260,
// 16'h5d55, 16'h566c, 16'h4db9, 16'h437f,
// 16'h37d9, 16'h2b20, 16'h1d7a, 16'h0f43,
// 16'h20bc, 16'hf22d, 16'he3eb, 16'hd639,
// 16'hc95b, 16'hbda1, 16'hb339, 16'haa5f,
// 16'ha349, 16'h9e07, 16'h9ad0, 16'h9999,
// 16'h9a7d, 16'h9d6e, 16'ha25d, 16'ha933,
// 16'hb1cb, 16'hbbf7, 16'hc789, 16'hd438,
// 16'he1d5, 16'hf020, 16'hfe8e, 16'h0d17,
// 16'h1b61, 16'h2920, 16'h3601, 16'h41d5,
// 16'h4c4a, 16'h5538, 16'h5c6a, 16'h61c0,
// 16'h6513, 16'h6667, 16'h6596, 16'h62c8,
// 16'h5ded, 16'h572f, 16'h4eaf, 16'h4490,
// 16'h3917, 16'h2c6d, 16'h1ee2, 16'h10b3,
// 16'h0231, 16'hf3a0, 16'he553, 16'hd78e,
// 16'hca9a, 16'hbebe, 16'hb431, 16'hab31,
// 16'ha3e6, 16'h9e7b, 16'h9b07, 16'h99a2,
// 16'h9a4f, 16'h9d0a, 16'ha1ca, 16'ha86c,
// 16'hb0df, 16'hbae1, 16'hc651, 16'hd2eb,
// 16'he06b, 16'hee96, 16'hfd15, 16'h0ba3,
// 16'h19fd, 16'h27c4, 16'h34c6, 16'h40b3,
// 16'h4b4e, 16'h546a, 16'h5bc5, 16'h614d,
// 16'h64d9, 16'h6656, 16'h65cb, 16'h6320,
// 16'h5e85, 16'h57ec, 16'h4f9f, 16'h45a3,
// 16'h3a4b, 16'h2dbd, 16'h2043, 16'h1226,
// 16'h03a4, 16'hf515, 16'he6bb, 16'hd8e6,
// 16'hcbdb, 16'hbfdf, 16'hb52e, 16'hac05,
// 16'ha48b, 16'h9eef, 16'h9b49, 16'h99ad,
// 16'h9a27, 16'h9cab, 16'ha13b, 16'ha7ae,
// 16'haff2, 16'hb9d0, 16'hc51f, 16'hd19b,
// 16'hdf0b, 16'hed25, 16'hfb9e, 16'h0a35,
// 16'h188d, 16'h266e, 16'h3384, 16'h3f8f,
// 16'h4a52, 16'h5390, 16'h5b1f, 16'h60d6,
// 16'h6494, 16'h664c, 16'h65eb, 16'h6382,
// 16'h5f0a, 16'h58b3, 16'h507f, 16'h46ba,
// 16'h3b78, 16'h2f0b, 16'h21a7, 16'h1392,
// 16'h051b, 16'hf689, 16'he824, 16'hda42,
// 16'hcd1c, 16'hc105, 16'hb62e, 16'hacde,
// 16'ha535, 16'h9f68, 16'h9b90, 16'h99bd,
// 16'h9a04, 16'h9c53, 16'ha0ae, 16'ha6f6,
// 16'haf09, 16'hb8c4, 16'hc3ed, 16'hd04f,
// 16'hddac, 16'hebb5, 16'hfa2a, 16'h08c1,
// 16'h1720, 16'h2517, 16'h323b, 16'h3e6e,
// 16'h4949, 16'h52bb, 16'h5a71, 16'h6059,
// 16'h644d, 16'h6635, 16'h6610, 16'h63d4,
// 16'h5f97, 16'h5965, 16'h516a, 16'h47c2,
// 16'h3ca9, 16'h3054, 16'h2307, 16'h14ff,
// 16'h0693, 16'hf7f9, 16'he993, 16'hdb9c,
// 16'hce62, 16'hc22d, 16'hb734, 16'hadb8,
// 16'ha5e6, 16'h9fe6, 16'h9bda, 16'h99d6,
// 16'h99e3, 16'h9c01, 16'ha02a, 16'ha63c,
// 16'hae29, 16'hb7b8, 16'hc2c0, 16'hcf09,
// 16'hdc49, 16'hea49, 16'hf8b5, 16'h074c,
// 16'h15b5, 16'h23b8, 16'h30f6, 16'h3d42,
// 16'h4846, 16'h51d9, 16'h59c1, 16'h5fd8,
// 16'h63fe, 16'h661f, 16'h6627, 16'h6429,
// 16'h6017, 16'h5a1c, 16'h5248, 16'h48cb,
// 16'h3dd3, 16'h319f, 16'h2462, 16'h1670,
// 16'h0804, 16'hf96e, 16'heb02, 16'hdcf7,
// 16'hcfae, 16'hc356, 16'hb83c, 16'hae9a,
// 16'ha697, 16'ha06d, 16'h9c28, 16'h99f4,
// 16'h99c7, 16'h9bb6, 16'h9fa6, 16'ha58e,
// 16'had48, 16'hb6b3, 16'hc197, 16'hcdbf,
// 16'hdaf1, 16'he8d8, 16'hf745, 16'h05d2,
// 16'h144d, 16'h2254, 16'h2fb2, 16'h3c11,
// 16'h473d, 16'h50f6, 16'h590b, 16'h5f53,
// 16'h63aa, 16'h6620, 16'h663e, 16'h6476,
// 16'h6092, 16'h5acf, 16'h5320, 16'h49d4,
// 16'h3efa, 16'h32e3, 16'h25c0, 16'h17d9,
// 16'h097a, 16'hfae5, 16'hec6c, 16'hde5b,
// 16'hd0f4, 16'hc487, 16'hb94a, 16'haf7c,
// 16'ha752, 16'ha0f3, 16'h9c80, 16'h9a13,
// 16'h99b5, 16'h9b6d, 16'h9f29, 16'ha4e3,
// 16'hac6c, 16'hb5b1, 16'hc070, 16'hcc7d,
// 16'hd991, 16'he773, 16'hf5cb, 16'h0462,
// 16'h12dc, 16'h20f3, 16'h2e68, 16'h3adf,
// 16'h4630, 16'h500f, 16'h5850, 16'h5ec9,
// 16'h6351, 16'h65dc, 16'h6651, 16'h64b8,
// 16'h6111, 16'h5b73, 16'h53fe, 16'h4ad0,
// 16'h4022, 16'h3425, 16'h2718, 16'h1948,
// 16'h0ae8, 16'hfc5f, 16'hedd8, 16'hdfbe,
// 16'hd242, 16'hc5b7, 16'hba5a, 16'hb065,
// 16'ha80f, 16'ha180, 16'h9cdc, 16'h9a38,
// 16'h99a9, 16'h9b26, 16'h9eb4, 16'ha43a,
// 16'hab97, 16'hb4b2, 16'hbf4d, 16'hcb3a,
// 16'hd83a, 16'he607, 16'hf459, 16'h02ed,
// 16'h116b, 16'h1f93, 16'h2d17, 16'h39ad,
// 16'h4520, 16'h4f22, 16'h5792, 16'h5e38,
// 16'h62f3, 16'h65b5, 16'h665b, 16'h64fa,
// 16'h6185, 16'h5c1a, 16'h54d0, 16'h4bcc,
// 16'h4146, 16'h3562, 16'h2875, 16'h1aad,
// 16'h0c5e, 16'hfdd1, 16'hef4b, 16'he120,
// 16'hd391, 16'hc6ed, 16'hbb6c, 16'hb153,
// 16'ha8d1, 16'ha211, 16'h9d3d, 16'h9a64,
// 16'h999e, 16'h9ae9, 16'h9e43, 16'ha394,
// 16'haaca, 16'hb3b3, 16'hbe2f, 16'hc9fa,
// 16'hd6e6, 16'he49a, 16'hf2ec, 16'h0170,
// 16'h1001, 16'h1e2b, 16'h2bc8, 16'h3877,
// 16'h4409, 16'h4e34, 16'h56cf, 16'h5da1,
// 16'h6293, 16'h6583, 16'h6666, 16'h6532,
// 16'h61f7, 16'h5cb9, 16'h559f, 16'h4cc8,
// 16'h4260, 16'h36a3, 16'h29c8, 16'h1c16,
// 16'h0dd2, 16'hff43, 16'hf0c0, 16'he281,
// 16'hd4e6, 16'hc822, 16'hbc84, 16'hb244,
// 16'ha997, 16'ha2a9, 16'h9da1, 16'h9a96,
// 16'h9998, 16'h9ab4, 16'h9dd1, 16'ha2fb,
// 16'ha9f8, 16'hb2bf, 16'hbd12, 16'hc8bf,
// 16'hd58e, 16'he337, 16'hf175, 16'h2020,
// 16'h0e8c, 16'h1cc7, 16'h2a74, 16'h373f,
// 16'h42f0, 16'h4d41, 16'h5606, 16'h5d08,
// 16'h622a, 16'h6552, 16'h6663, 16'h656d,
// 16'h625e, 16'h5d56, 16'h566b, 16'h4dbb,
// 16'h437b, 16'h37e0, 16'h2b18, 16'h1d81,
// 16'h0f3f, 16'h20bd, 16'hf22e, 16'he3ea,
// 16'hd638, 16'hc95e, 16'hbd9e, 16'hb33a,
// 16'haa60, 16'ha346, 16'h9e0c, 16'h9aca,
// 16'h999e, 16'h9a7a, 16'h9d70, 16'ha25c,
// 16'ha933, 16'hb1cb, 16'hbbf8, 16'hc787,
// 16'hd43c, 16'he1d0, 16'hf004, 16'hfe8c,
// 16'h0d16, 16'h1b64, 16'h291d, 16'h3605,
// 16'h41d1, 16'h4c4c, 16'h5537, 16'h5c6b,
// 16'h61bf, 16'h6515, 16'h6664, 16'h6599,
// 16'h62c6, 16'h5ded, 16'h5730, 16'h4ead,
// 16'h4493, 16'h3914, 16'h2c6f, 16'h1ee0,
// 16'h10b4, 16'h0230, 16'hf3a2, 16'he551,
// 16'hd78f, 16'hca9a, 16'hbebc, 16'hb435,
// 16'hab2d, 16'ha3e9, 16'h9e78, 16'h9b09,
// 16'h99a2, 16'h9a4e, 16'h9d0c, 16'ha1c6,
// 16'ha871, 16'hb0da, 16'hbae4, 16'hc651,
// 16'hd2e9, 16'he06f, 16'hee92, 16'hfd16,
// 16'h0ba5, 16'h19f9, 16'h27c8, 16'h34c4,
// 16'h40b5, 16'h4b4c, 16'h546a, 16'h5bc5,
// 16'h614e, 16'h64d8, 16'h6657, 16'h65c9,
// 16'h6323, 16'h5e82, 16'h57ef, 16'h4f9c,
// 16'h45a5, 16'h3a4a, 16'h2dbd, 16'h2044,
// 16'h1224, 16'h03a6, 16'hf515, 16'he6b9,
// 16'hd8e8, 16'hcbd8, 16'hbfe2, 16'hb52d,
// 16'hac05, 16'ha48b, 16'h9eef, 16'h9b48,
// 16'h99af, 16'h9a24, 16'h9cb0, 16'ha136,
// 16'ha7b1, 16'haff0, 16'hb9d1, 16'hc51f,
// 16'hd19c, 16'hdf0a, 16'hed25, 16'hfb9e,
// 16'h0a34, 16'h188f, 16'h266d, 16'h3385,
// 16'h3f8e, 16'h4a52, 16'h5391, 16'h5b1e,
// 16'h60d7, 16'h6493, 16'h664c, 16'h65ec,
// 16'h6380, 16'h5f0d, 16'h58af, 16'h5082,
// 16'h46b8, 16'h3b79, 16'h2f0b, 16'h21a6,
// 16'h1393, 16'h051b, 16'hf688, 16'he825,
// 16'hda41, 16'hcd1d, 16'hc104, 16'hb630,
// 16'hacdb, 16'ha537, 16'h9f68, 16'h9b8e,
// 16'h99c1, 16'h99ff, 16'h9c57, 16'ha0ad,
// 16'ha6f5, 16'haf09, 16'hb8c5, 16'hc3eb,
// 16'hd053, 16'hdda8, 16'hebb6, 16'hfa2c,
// 16'h08bc, 16'h1726, 16'h2512, 16'h323f,
// 16'h3e6a, 16'h494d, 16'h52b7, 16'h5a74,
// 16'h6057, 16'h644e, 16'h6635, 16'h6610,
// 16'h63d4, 16'h5f96, 16'h5967, 16'h5167,
// 16'h47c5, 16'h3ca6, 16'h3057, 16'h2305,
// 16'h1520, 16'h0692, 16'hf7f9, 16'he995,
// 16'hdb9a, 16'hce63, 16'hc22d, 16'hb733,
// 16'hadba, 16'ha5e3, 16'h9fe9, 16'h9bd8,
// 16'h99d8, 16'h99e1, 16'h9c03, 16'ha027,
// 16'ha640, 16'hae26, 16'hb7b9, 16'hc2c2,
// 16'hcf04, 16'hdc4f, 16'hea44, 16'hf8ba,
// 16'h0747, 16'h15b9, 16'h23b5, 16'h30f9,
// 16'h3d40, 16'h4846, 16'h51d9, 16'h59c2,
// 16'h5fd7, 16'h63ff, 16'h661d, 16'h6629,
// 16'h6428, 16'h6017, 16'h5a1c, 16'h5248,
// 16'h48ca, 16'h3dd7, 16'h319a, 16'h2466,
// 16'h166d, 16'h0805, 16'hf970, 16'heafe,
// 16'hdcfd, 16'hcfa6, 16'hc35e, 16'hb837,
// 16'hae9c, 16'ha698, 16'ha069, 16'h9c2d,
// 16'h99f0, 16'h99ca, 16'h9bb4, 16'h9fa7,
// 16'ha58d, 16'had49, 16'hb6b2, 16'hc197,
// 16'hcdc1, 16'hdaed, 16'he8dd, 16'hf740,
// 16'h05d6, 16'h144a, 16'h2257, 16'h2faf,
// 16'h3c13, 16'h473c, 16'h50f7, 16'h590a,
// 16'h5f53, 16'h63aa, 16'h6601, 16'h663e,
// 16'h6474, 16'h6094, 16'h5acd, 16'h5322,
// 16'h49d2, 16'h3efb, 16'h32e4, 16'h25be,
// 16'h17db, 16'h0977, 16'hfae7, 16'hec6c,
// 16'hde5b, 16'hd0f4, 16'hc486, 16'hb94b,
// 16'haf7a, 16'ha755, 16'ha0f0, 16'h9c81,
// 16'h9a15, 16'h99b2, 16'h9b6f, 16'h9f27,
// 16'ha4e4, 16'hac6d, 16'hb5af, 16'hc072,
// 16'hcc7a, 16'hd995, 16'he76f, 16'hf5cf,
// 16'h045e, 16'h12de, 16'h20f4, 16'h2e65,
// 16'h3ae2, 16'h462e, 16'h5010, 16'h5851,
// 16'h5ec6, 16'h6353, 16'h65da, 16'h6654,
// 16'h64b5, 16'h6113, 16'h5b74, 16'h53fa,
// 16'h4ad5, 16'h401c, 16'h342a, 16'h2717,
// 16'h1946, 16'h0aec, 16'hfc59, 16'heddd,
// 16'hdfbc, 16'hd241, 16'hc5ba, 16'hba56,
// 16'hb068, 16'ha80e, 16'ha180, 16'h9cdc,
// 16'h9a39, 16'h99a7, 16'h9b28, 16'h9eb4,
// 16'ha437, 16'hab9c, 16'hb4ae, 16'hbf4f,
// 16'hcb3a, 16'hd838, 16'he609, 16'hf458,
// 16'h02ed, 16'h116a, 16'h1f95, 16'h2d14,
// 16'h39b1, 16'h451b, 16'h4f26, 16'h5790,
// 16'h5e37, 16'h62f7, 16'h65b0, 16'h665f,
// 16'h64f8, 16'h6185, 16'h5c1a, 16'h54d1,
// 16'h4bcb, 16'h4147, 16'h3561, 16'h2875,
// 16'h1aad, 16'h0c5e, 16'hfdd2, 16'hef49,
// 16'he122, 16'hd390, 16'hc6ec, 16'hbb6e,
// 16'hb152, 16'ha8d0, 16'ha214, 16'h9d39,
// 16'h9a68, 16'h999b, 16'h9aec, 16'h9e40,
// 16'ha397, 16'haac6, 16'hb3b7, 16'hbe2d,
// 16'hc9fc, 16'hd6e2, 16'he49f, 16'hf2e6,
// 16'h0177, 16'h0ffb, 16'h1e2f, 16'h2bc6,
// 16'h3878, 16'h4408, 16'h4e34, 16'h56d0,
// 16'h5d9f, 16'h6296, 16'h6581, 16'h6665,
// 16'h6535, 16'h61f3, 16'h5cbc, 16'h559f,
// 16'h4cc6, 16'h4262, 16'h36a2, 16'h29c8,
// 16'h1c17, 16'h0dd0, 16'hff46, 16'hf0bc,
// 16'he285, 16'hd4e3, 16'hc823, 16'hbc85,
// 16'hb243, 16'ha997, 16'ha2a9, 16'h9da2,
// 16'h9a93, 16'h999e, 16'h9aad, 16'h9dd7,
// 16'ha2f6, 16'ha9fc, 16'hb2bc, 16'hbd14,
// 16'hc8be, 16'hd58e, 16'he336, 16'hf177,
// 16'hfffe, 16'h0e8d, 16'h1cc7, 16'h2a74,
// 16'h373f, 16'h42ef, 16'h4d42, 16'h5605,
// 16'h5d0a, 16'h6229, 16'h6551, 16'h6665,
// 16'h656b, 16'h625f, 16'h5d56, 16'h566b,
// 16'h4dbb, 16'h437c, 16'h37dd, 16'h2b1c,
// 16'h1d7c, 16'h0f44, 16'h20ba, 16'hf22f,
// 16'he3ea, 16'hd637, 16'hc95e, 16'hbda0,
// 16'hb338, 16'haa61, 16'ha345, 16'h9e0c,
// 16'h9acc, 16'h999c, 16'h9a7c, 16'h9d6d,
// 16'ha25e, 16'ha932, 16'hb1cb, 16'hbbf9,
// 16'hc787, 16'hd43a, 16'he1d1, 16'hf005,
// 16'hfe8a, 16'h0d19, 16'h1b62, 16'h291d,
// 16'h3605, 16'h41d2, 16'h4c4b, 16'h5537,
// 16'h5c6c, 16'h61be, 16'h6515, 16'h6665,
// 16'h6596, 16'h62ca, 16'h5de9, 16'h5733,
// 16'h4eab, 16'h4494, 16'h3914, 16'h2c6f,
// 16'h1edf, 16'h10b6, 16'h022e, 16'hf3a3,
// 16'he552, 16'hd78d, 16'hca9b, 16'hbebd,
// 16'hb433, 16'hab2e, 16'ha3ea, 16'h9e76,
// 16'h9b0c, 16'h999f, 16'h9a4f, 16'h9d0c,
// 16'ha1c7, 16'ha871, 16'hb0d9, 16'hbae5,
// 16'hc64f, 16'hd2ec, 16'he06b, 16'hee96,
// 16'hfd13, 16'h0ba7, 16'h19f9, 16'h27c6,
// 16'h34c6, 16'h40b2, 16'h4b50, 16'h5467,
// 16'h5bc7, 16'h614d, 16'h64d7, 16'h665a,
// 16'h65c6, 16'h6324, 16'h5e82, 16'h57ef,
// 16'h4f9c, 16'h45a6, 16'h3a49, 16'h2dbd,
// 16'h2045, 16'h1223, 16'h03a7, 16'hf513,
// 16'he6bc, 16'hd8e5, 16'hcbdb, 16'hbfe0,
// 16'hb52e, 16'hac04, 16'ha48c, 16'h9eee,
// 16'h9b4a, 16'h99ad, 16'h9a26, 16'h9cad,
// 16'ha139, 16'ha7ae, 16'haff3, 16'hb9cf,
// 16'hc521, 16'hd199, 16'hdf0b, 16'hed26,
// 16'hfb9d, 16'h0a36, 16'h188c, 16'h266f,
// 16'h3384, 16'h3f8e, 16'h4a53, 16'h538e,
// 16'h5b23, 16'h60d2, 16'h6496, 16'h664b,
// 16'h65eb, 16'h6383, 16'h5f0a, 16'h58b1,
// 16'h5081, 16'h46b8, 16'h3b7a, 16'h2f0a,
// 16'h21a7, 16'h1391, 16'h051d, 16'hf685,
// 16'he829, 16'hda3d, 16'hcd20, 16'hc102,
// 16'hb630, 16'hacdd, 16'ha534, 16'h9f6b,
// 16'h9b8c, 16'h99c1, 16'h9a01, 16'h9c55,
// 16'ha0ad, 16'ha6f6, 16'haf08, 16'hb8c6,
// 16'hc3ec, 16'hd051, 16'hdda8, 16'hebb8,
// 16'hfa28, 16'h08c3, 16'h171e, 16'h2518,
// 16'h323b, 16'h3e6d, 16'h494b, 16'h52b9,
// 16'h5a71, 16'h605a, 16'h644c, 16'h6636,
// 16'h6610, 16'h63d3, 16'h5f98, 16'h5964,
// 16'h516b, 16'h47c0, 16'h3cab, 16'h3054,
// 16'h2305, 16'h1504, 16'h068c, 16'hf7ff,
// 16'he98f, 16'hdb9f, 16'hce61, 16'hc22d,
// 16'hb734, 16'hadb8, 16'ha5e6, 16'h9fe5,
// 16'h9bdc, 16'h99d4, 16'h99e5, 16'h9c01,
// 16'ha027, 16'ha640, 16'hae26, 16'hb7b9,
// 16'hc2c2, 16'hcf06, 16'hdc4b, 16'hea49,
// 16'hf8b4, 16'h074c, 16'h15b7, 16'h23b5,
// 16'h30fa, 16'h3d3e, 16'h4849, 16'h51d7,
// 16'h59c2, 16'h5fd8, 16'h63fe, 16'h661e,
// 16'h6629, 16'h6428, 16'h6016, 16'h5a1e,
// 16'h5245, 16'h48cd, 16'h3dd5, 16'h319b,
// 16'h2466, 16'h166c, 16'h0806, 16'hf96e,
// 16'heb02, 16'hdcf8, 16'hcfac, 16'hc357,
// 16'hb83d, 16'hae98, 16'ha69b, 16'ha068,
// 16'h9c2c, 16'h99f2, 16'h99c8, 16'h9bb7,
// 16'h9fa3, 16'ha591, 16'had46, 16'hb6b4,
// 16'hc196, 16'hcdc2, 16'hdaeb, 16'he8de,
// 16'hf740, 16'h05d6, 16'h144b, 16'h2256,
// 16'h2fae, 16'h3c15, 16'h473a, 16'h50f9,
// 16'h590a, 16'h5f51, 16'h63ad, 16'h65fd,
// 16'h6642, 16'h6471, 16'h6097, 16'h5aca,
// 16'h5324, 16'h49d1, 16'h3efb, 16'h32e5,
// 16'h25bd, 16'h17db, 16'h0979, 16'hfae4,
// 16'hec6e, 16'hde5a, 16'hd0f5, 16'hc487,
// 16'hb948, 16'haf7e, 16'ha750, 16'ha0f4,
// 16'h9c81, 16'h9a11, 16'h99b8, 16'h9b6a,
// 16'h9f2a, 16'ha4e2, 16'hac6e, 16'hb5b0,
// 16'hc071, 16'hcc7c, 16'hd990, 16'he774,
// 16'hf5cb, 16'h0464, 16'h12d7, 16'h20f9,
// 16'h2e62, 16'h3ae3, 16'h462f, 16'h500e,
// 16'h5852, 16'h5ec6, 16'h6354, 16'h65d9,
// 16'h6654, 16'h64b6, 16'h6111, 16'h5b75,
// 16'h53fb, 16'h4ad3, 16'h401f, 16'h3427,
// 16'h2719, 16'h1945, 16'h0aec, 16'hfc5a,
// 16'heddc, 16'hdfbc, 16'hd242, 16'hc5b9,
// 16'hba57, 16'hb067, 16'ha80e, 16'ha181,
// 16'h9cdb, 16'h9a3a, 16'h99a4, 16'h9b2c,
// 16'h9eb0, 16'ha43c, 16'hab97, 16'hb4b1,
// 16'hbf4d, 16'hcb3b, 16'hd839, 16'he608,
// 16'hf459, 16'h02ec, 16'h116b, 16'h1f93,
// 16'h2d17, 16'h39ae, 16'h451e, 16'h4f23,
// 16'h5792, 16'h5e37, 16'h62f5, 16'h65b2,
// 16'h665e, 16'h64f7, 16'h6188, 16'h5c17,
// 16'h54d2, 16'h4bcd, 16'h4142, 16'h3567,
// 16'h2871, 16'h1aae, 16'h0c61, 16'hfdcc,
// 16'hef50, 16'he11b, 16'hd396, 16'hc6e9,
// 16'hbb6e, 16'hb153, 16'ha8cf, 16'ha214,
// 16'h9d3b, 16'h9a64, 16'h999f, 16'h9ae9,
// 16'h9e42, 16'ha396, 16'haac7, 16'hb3b5,
// 16'hbe2f, 16'hc9fb, 16'hd6e2, 16'he49f,
// 16'hf2e6, 16'h0177, 16'h0ffc, 16'h1e2d,
// 16'h2bc8, 16'h3876, 16'h440b, 16'h4e32,
// 16'h56d0, 16'h5da1, 16'h6293, 16'h6584,
// 16'h6664, 16'h6534, 16'h61f5, 16'h5cb9,
// 16'h55a2, 16'h4cc4, 16'h4263, 16'h36a2,
// 16'h29c7, 16'h1c18, 16'h0dcf, 16'hff47,
// 16'hf0bc, 16'he284, 16'hd4e4, 16'hc823,
// 16'hbc84, 16'hb245, 16'ha994, 16'ha2ac,
// 16'h9d9f, 16'h9a96, 16'h999c, 16'h9aad,
// 16'h9dd8, 16'ha2f5, 16'ha9fc, 16'hb2bf,
// 16'hbd0f, 16'hc8c2, 16'hd58b, 16'he33a,
// 16'hf173, 16'h2001, 16'h0e8a, 16'h1cc9,
// 16'h2a74, 16'h373e, 16'h42f0, 16'h4d41,
// 16'h5606, 16'h5d09, 16'h622a, 16'h6550,
// 16'h6667, 16'h6568, 16'h6262, 16'h5d54,
// 16'h566b, 16'h4dbc, 16'h437b, 16'h37dd,
// 16'h2b1d, 16'h1d7c, 16'h0f42, 16'h20bd,
// 16'hf22c, 16'he3ec, 16'hd638, 16'hc95c,
// 16'hbda0, 16'hb339, 16'haa60, 16'ha348,
// 16'h9e09, 16'h9acd, 16'h999a, 16'h9a7f,
// 16'h9d6c, 16'ha25f, 16'ha930, 16'hb1cd,
// 16'hbbf7, 16'hc788, 16'hd43b, 16'he1d0,
// 16'hf004, 16'hfe8d, 16'h0d15, 16'h1b65,
// 16'h291c, 16'h3604, 16'h41d3, 16'h4c4b,
// 16'h5538, 16'h5c6b, 16'h61bd, 16'h6517,
// 16'h6662, 16'h659c, 16'h62c4, 16'h5ded,
// 16'h5731, 16'h4eac, 16'h4494, 16'h3913,
// 16'h2c70, 16'h1edf, 16'h10b6, 16'h022e,
// 16'hf3a2, 16'he553, 16'hd78c, 16'hca9c,
// 16'hbebd, 16'hb431, 16'hab31, 16'ha3e7,
// 16'h9e78, 16'h9b0b, 16'h999f, 16'h9a50,
// 16'h9d0b, 16'ha1c7, 16'ha871, 16'hb0da,
// 16'hbae3, 16'hc652, 16'hd2e9, 16'he06e,
// 16'hee93, 16'hfd16, 16'h0ba4, 16'h19fc,
// 16'h27c3, 16'h34c8, 16'h40b1, 16'h4b51,
// 16'h5466, 16'h5bc8, 16'h614a, 16'h64dc,
// 16'h6655, 16'h65ca, 16'h6322, 16'h5e81,
// 16'h57f3, 16'h4f98, 16'h45a8, 16'h3a48,
// 16'h2dbe, 16'h2044, 16'h1225, 16'h03a4,
// 16'hf515, 16'he6bb, 16'hd8e6, 16'hcbdc,
// 16'hbfdd, 16'hb530, 16'hac02, 16'ha48e,
// 16'h9eee, 16'h9b49, 16'h99ae, 16'h9a23,
// 16'h9cb0, 16'ha137, 16'ha7b1, 16'haff0,
// 16'hb9d1, 16'hc51e, 16'hd19c, 16'hdf0a,
// 16'hed26, 16'hfb9e, 16'h0a33, 16'h1890,
// 16'h266c, 16'h3386, 16'h3f8d, 16'h4a53,
// 16'h538f, 16'h5b22, 16'h60d3, 16'h6495,
// 16'h664c, 16'h65ea, 16'h6384, 16'h5f09,
// 16'h58b1, 16'h5082, 16'h46b7, 16'h3b7b,
// 16'h2f09, 16'h21a6, 16'h1394, 16'h051b,
// 16'hf686, 16'he829, 16'hda3c, 16'hcd22,
// 16'hc120, 16'hb633, 16'hacda, 16'ha537,
// 16'h9f68, 16'h9b8e, 16'h99c2, 16'h99fe,
// 16'h9c58, 16'ha0ac, 16'ha6f4, 16'haf0d,
// 16'hb8c0, 16'hc3f0, 16'hd04f, 16'hdda9,
// 16'hebb7, 16'hfa2a, 16'h08c0, 16'h1722,
// 16'h2513, 16'h323f, 16'h3e6a, 16'h494e,
// 16'h52b7, 16'h5a72, 16'h6059, 16'h644d,
// 16'h6636, 16'h660e, 16'h63d6, 16'h5f95,
// 16'h5967, 16'h5169, 16'h47c1, 16'h3ca9,
// 16'h3056, 16'h2304, 16'h1503, 16'h068f,
// 16'hf7fc, 16'he992, 16'hdb9c, 16'hce63,
// 16'hc22b, 16'hb737, 16'hadb6, 16'ha5e7,
// 16'h9fe4, 16'h9bde, 16'h99d2, 16'h99e6,
// 16'h9c20, 16'ha028, 16'ha63f, 16'hae27,
// 16'hb7b9, 16'hc2c1, 16'hcf07, 16'hdc4a,
// 16'hea49, 16'hf8b4, 16'h074e, 16'h15b2,
// 16'h23bb, 16'h30f5, 16'h3d41, 16'h4847,
// 16'h51d8, 16'h59c1, 16'h5fda, 16'h63fc,
// 16'h661f, 16'h6629, 16'h6426, 16'h601a,
// 16'h5a19, 16'h524a, 16'h48ca, 16'h3dd5,
// 16'h319d, 16'h2462, 16'h1671, 16'h0801,
// 16'hf974, 16'heafc, 16'hdcfb, 16'hcfac,
// 16'hc356, 16'hb83e, 16'hae98, 16'ha699,
// 16'ha06b, 16'h9c2a, 16'h99f2, 16'h99c9,
// 16'h9bb5, 16'h9fa6, 16'ha58e, 16'had48,
// 16'hb6b3, 16'hc196, 16'hcdc2, 16'hdaec,
// 16'he8dd, 16'hf741, 16'h05d5, 16'h144c,
// 16'h2254, 16'h2fb1, 16'h3c13, 16'h473a,
// 16'h50fa, 16'h5908, 16'h5f54, 16'h63ab,
// 16'h65fd, 16'h6643, 16'h646f, 16'h609a,
// 16'h5ac7, 16'h5328, 16'h49cc, 16'h3f20,
// 16'h32df, 16'h25c3, 16'h17d8, 16'h097a,
// 16'hfae3, 16'hec6f, 16'hde59, 16'hd0f6,
// 16'hc486, 16'hb948, 16'haf7f, 16'ha750,
// 16'ha0f4, 16'h9c80, 16'h9a12, 16'h99b7,
// 16'h9b6a, 16'h9f2c, 16'ha4e0, 16'hac6f,
// 16'hb5b0, 16'hc070, 16'hcc7c, 16'hd993,
// 16'he76f, 16'hf5d0, 16'h045f, 16'h12dc,
// 16'h20f6, 16'h2e63, 16'h3ae3, 16'h462e,
// 16'h5010, 16'h5850, 16'h5ec8, 16'h6353,
// 16'h65d8, 16'h6656, 16'h64b3, 16'h6116,
// 16'h5b70, 16'h53fe, 16'h4ad1, 16'h4020,
// 16'h3427, 16'h2718, 16'h1947, 16'h0aea,
// 16'hfc5c, 16'hedda, 16'hdfbe, 16'hd240,
// 16'hc5bb, 16'hba55, 16'hb06a, 16'ha80c,
// 16'ha180, 16'h9cdd, 16'h9a37, 16'h99a9,
// 16'h9b27, 16'h9eb4, 16'ha438, 16'hab9a,
// 16'hb4af, 16'hbf50, 16'hcb38, 16'hd83b,
// 16'he606, 16'hf45a, 16'h02ee, 16'h1168,
// 16'h1f96, 16'h2d13, 16'h39b2, 16'h451b,
// 16'h4f26, 16'h578f, 16'h5e39, 16'h62f4,
// 16'h65b2, 16'h665f, 16'h64f7, 16'h6187,
// 16'h5c18, 16'h54d1, 16'h4bcd, 16'h4144,
// 16'h3565, 16'h2871, 16'h1aaf, 16'h0c5e,
// 16'hfdd0, 16'hef4d, 16'he11d, 16'hd394,
// 16'hc6ea, 16'hbb6e, 16'hb152, 16'ha8d2,
// 16'ha210, 16'h9d3e, 16'h9a63, 16'h999e,
// 16'h9aec, 16'h9e3e, 16'ha39a, 16'haac3,
// 16'hb3b9, 16'hbe2b, 16'hc9fe, 16'hd6e1,
// 16'he49f, 16'hf2e6, 16'h0178, 16'h0ff8,
// 16'h1e32, 16'h2bc4, 16'h3879, 16'h4409,
// 16'h4e33, 16'h56ce, 16'h5da3, 16'h6292,
// 16'h6584, 16'h6664, 16'h6535, 16'h61f2,
// 16'h5cbf, 16'h559a, 16'h4ccb, 16'h425f,
// 16'h36a3, 16'h29c9, 16'h1c14, 16'h0dd3,
// 16'hff44, 16'hf0be, 16'he284, 16'hd4e3,
// 16'hc823, 16'hbc85, 16'hb243, 16'ha998,
// 16'ha2a8, 16'h9da2, 16'h9a94, 16'h999c,
// 16'h9aaf, 16'h9dd7, 16'ha2f4, 16'ha9fe,
// 16'hb2bb, 16'hbd15, 16'hc8bc, 16'hd591,
// 16'he333, 16'hf178, 16'h2020, 16'h0e89,
// 16'h1ccb, 16'h2a71, 16'h3741, 16'h42ee,
// 16'h4d43, 16'h5603, 16'h5d0c, 16'h6228,
// 16'h6552, 16'h6664, 16'h656b, 16'h625e,
// 16'h5d59, 16'h5667, 16'h4dbe, 16'h437b,
// 16'h37dc, 16'h2b1e, 16'h1d7b, 16'h0f43,
// 16'h20bc, 16'hf22d, 16'he3ec, 16'hd637,
// 16'hc95c, 16'hbda2, 16'hb336, 16'haa64,
// 16'ha343, 16'h9e0c, 16'h9acb, 16'h999f,
// 16'h9a77, 16'h9d74, 16'ha257, 16'ha938,
// 16'hb1c7, 16'hbbfb, 16'hc785, 16'hd43d,
// 16'he1cf, 16'hf006, 16'hfe89, 16'h0d19,
// 16'h1b63, 16'h291b, 16'h3608, 16'h41cd,
// 16'h4c51, 16'h5533, 16'h5c6e, 16'h61bc,
// 16'h6516, 16'h6665, 16'h6597, 16'h62c9,
// 16'h5dea, 16'h5732, 16'h4eac, 16'h4493,
// 16'h3915, 16'h2c6d, 16'h1ee2, 16'h10b3,
// 16'h0231, 16'hf3a2, 16'he550, 16'hd78f,
// 16'hca9a, 16'hbebd, 16'hb433, 16'hab2f,
// 16'ha3e9, 16'h9e76, 16'h9b0c, 16'h999e,
// 16'h9a52, 16'h9d08, 16'ha1ca, 16'ha86e,
// 16'hb0dd, 16'hbae2, 16'hc651, 16'hd2ea,
// 16'he06d, 16'hee95, 16'hfd13, 16'h0ba8,
// 16'h19f6, 16'h27cb, 16'h34c1, 16'h40b6,
// 16'h4b4e, 16'h5466, 16'h5bca, 16'h6149,
// 16'h64db, 16'h6657, 16'h65c8, 16'h6323,
// 16'h5e82, 16'h57ef, 16'h4f9c, 16'h45a6,
// 16'h3a49, 16'h2dbd, 16'h2045, 16'h1223,
// 16'h03a7, 16'hf512, 16'he6be, 16'hd8e4,
// 16'hcbdc, 16'hbfde, 16'hb52f, 16'hac03,
// 16'ha48e, 16'h9eed, 16'h9b4a, 16'h99ae,
// 16'h9a23, 16'h9cb0, 16'ha136, 16'ha7b3,
// 16'hafee, 16'hb9d3, 16'hc51c, 16'hd19d,
// 16'hdf0a, 16'hed25, 16'hfb9f, 16'h0a34,
// 16'h188c, 16'h2671, 16'h3381, 16'h3f92,
// 16'h4a4f, 16'h5392, 16'h5b1e, 16'h60d6,
// 16'h6495, 16'h664a, 16'h65ee, 16'h637e,
// 16'h5f0e, 16'h58ae, 16'h5084, 16'h46b6,
// 16'h3b7a, 16'h2f0b, 16'h21a6, 16'h1393,
// 16'h051a, 16'hf689, 16'he824, 16'hda44,
// 16'hcd19, 16'hc108, 16'hb62c, 16'hacde,
// 16'ha536, 16'h9f67, 16'h9b92, 16'h99bb,
// 16'h9a05, 16'h9c52, 16'ha0af, 16'ha6f6,
// 16'haf08, 16'hb8c5, 16'hc3ec, 16'hd051,
// 16'hddaa, 16'hebb6, 16'hfa2a, 16'h08bf,
// 16'h1724, 16'h2513, 16'h323e, 16'h3e6b,
// 16'h494c, 16'h52b9, 16'h5a72, 16'h6059,
// 16'h644b, 16'h6639, 16'h660a, 16'h63da,
// 16'h5f92, 16'h596a, 16'h5166, 16'h47c3,
// 16'h3ca9, 16'h3054, 16'h2308, 16'h14ff,
// 16'h0691, 16'hf7fc, 16'he990, 16'hdb9f,
// 16'hce60, 16'hc22e, 16'hb733, 16'hadb9,
// 16'ha5e5, 16'h9fe7, 16'h9bda, 16'h99d5,
// 16'h99e3, 16'h9c03, 16'ha027, 16'ha63f,
// 16'hae27, 16'hb7b9, 16'hc2c0, 16'hcf08,
// 16'hdc4a, 16'hea49, 16'hf8b6, 16'h0749,
// 16'h15b9, 16'h23b4, 16'h30fa, 16'h3d3f,
// 16'h4847, 16'h51d9, 16'h59c2, 16'h5fd6,
// 16'h6420, 16'h661c, 16'h662c, 16'h6424,
// 16'h601b, 16'h5a18, 16'h524b, 16'h48ca,
// 16'h3dd4, 16'h319e, 16'h2462, 16'h1670,
// 16'h0803, 16'hf972, 16'heafd, 16'hdcfb,
// 16'hcfab, 16'hc357, 16'hb83e, 16'hae97,
// 16'ha69a, 16'ha06a, 16'h9c2b, 16'h99f1,
// 16'h99ca, 16'h9bb3, 16'h9fa9, 16'ha58b,
// 16'had4a, 16'hb6b2, 16'hc198, 16'hcdbe,
// 16'hdaf1, 16'he8d7, 16'hf746, 16'h05d4,
// 16'h144a, 16'h2256, 16'h2faf, 16'h3c14,
// 16'h473b, 16'h50f9, 16'h5907, 16'h5f56,
// 16'h63a9, 16'h65ff, 16'h6641, 16'h6471,
// 16'h6097, 16'h5acc, 16'h5322, 16'h49d2,
// 16'h3efb, 16'h32e3, 16'h25bf, 16'h17db,
// 16'h0978, 16'hfae5, 16'hec6e, 16'hde59,
// 16'hd0f6, 16'hc485, 16'hb94a, 16'haf7c,
// 16'ha754, 16'ha0f0, 16'h9c83, 16'h9a11,
// 16'h99b5, 16'h9b6e, 16'h9f28, 16'ha4e3,
// 16'hac6d, 16'hb5b0, 16'hc071, 16'hcc7b,
// 16'hd995, 16'he76d, 16'hf5d1, 16'h045e,
// 16'h12dd, 16'h20f5, 16'h2e64, 16'h3ae2,
// 16'h462f, 16'h5010, 16'h584f, 16'h5ec8,
// 16'h6353, 16'h65da, 16'h6653, 16'h64b6,
// 16'h6112, 16'h5b74, 16'h53fc, 16'h4ad1,
// 16'h4021, 16'h3426, 16'h2719, 16'h1946,
// 16'h0aeb, 16'hfc5a, 16'heddd, 16'hdfbb,
// 16'hd243, 16'hc5b8, 16'hba58, 16'hb066,
// 16'ha80f, 16'ha180, 16'h9cdc, 16'h9a38,
// 16'h99a8, 16'h9b27, 16'h9eb5, 16'ha438,
// 16'hab99, 16'hb4b1, 16'hbf4c, 16'hcb3d,
// 16'hd837, 16'he608, 16'hf45b, 16'h02e9,
// 16'h116e, 16'h1f91, 16'h2d18, 16'h39ae,
// 16'h451d, 16'h4f25, 16'h5790, 16'h5e39,
// 16'h62f4, 16'h65b1, 16'h6661, 16'h64f4,
// 16'h618b, 16'h5c14, 16'h54d4, 16'h4bcb,
// 16'h4145, 16'h3564, 16'h2873, 16'h1aad,
// 16'h0c60, 16'hfdcf, 16'hef4d, 16'he11e,
// 16'hd392, 16'hc6ec, 16'hbb6d, 16'hb153,
// 16'ha8d0, 16'ha212, 16'h9d3c, 16'h9a64,
// 16'h999f, 16'h9ae8, 16'h9e44, 16'ha393,
// 16'haacb, 16'hb3b2, 16'hbe31, 16'hc9f9,
// 16'hd6e4, 16'he49d, 16'hf2e9, 16'h0175,
// 16'h0ffb, 16'h1e30, 16'h2bc3, 16'h387d,
// 16'h4404, 16'h4e37, 16'h56cd, 16'h5da2,
// 16'h6293, 16'h6584, 16'h6663, 16'h6536,
// 16'h61f3, 16'h5cbc, 16'h559d, 16'h4cc9,
// 16'h425f, 16'h36a5, 16'h29c6, 16'h1c18,
// 16'h0dcf, 16'hff47, 16'hf0bd, 16'he282,
// 16'hd4e7, 16'hc820, 16'hbc87, 16'hb242,
// 16'ha998, 16'ha2a7, 16'h9da5, 16'h9a92,
// 16'h999c, 16'h9ab0, 16'h9dd5, 16'ha2f7,
// 16'ha9fb, 16'hb2be, 16'hbd11, 16'hc8c1,
// 16'hd58b, 16'he339, 16'hf175, 16'hffff,
// 16'h0e8d, 16'h1cc5, 16'h2a77, 16'h373d,
// 16'h42f1, 16'h4d41, 16'h5605, 16'h5d08,
// 16'h622d, 16'h654e, 16'h6668, 16'h6567,
// 16'h6262, 16'h5d54, 16'h566d, 16'h4db9,
// 16'h437d, 16'h37dc, 16'h2b1d, 16'h1d7c,
// 16'h0f43, 16'h20ba, 16'hf230, 16'he3e9,
// 16'hd639, 16'hc95c, 16'hbda0, 16'hb339,
// 16'haa61, 16'ha345, 16'h9e0c, 16'h9acc,
// 16'h999b, 16'h9a7d, 16'h9d6d, 16'ha25e,
// 16'ha932, 16'hb1cc, 16'hbbf7, 16'hc788,
// 16'hd43b, 16'he1cf, 16'hf007, 16'hfe88,
// 16'h0d1b, 16'h1b60, 16'h291e, 16'h3604,
// 16'h41d3, 16'h4c4a, 16'h553a, 16'h5c67,
// 16'h61c2, 16'h6513, 16'h6665, 16'h6599,
// 16'h62c6, 16'h5dec, 16'h5732, 16'h4eac,
// 16'h4492, 16'h3916, 16'h2c6c, 16'h1ee4,
// 16'h10b2, 16'h0231, 16'hf39f, 16'he555,
// 16'hd78b, 16'hca9d, 16'hbebc, 16'hb431,
// 16'hab32, 16'ha3e4, 16'h9e7d, 16'h9b05,
// 16'h99a5, 16'h9a4c, 16'h9d0d, 16'ha1c7,
// 16'ha86f, 16'hb0dc, 16'hbae4, 16'hc650,
// 16'hd2eb, 16'he06b, 16'hee96, 16'hfd14,
// 16'h0ba6, 16'h19f9, 16'h27c7, 16'h34c5,
// 16'h40b4, 16'h4b4e, 16'h5468, 16'h5bc6,
// 16'h614d, 16'h64d9, 16'h6658, 16'h65c8,
// 16'h6323, 16'h5e80, 16'h57f3, 16'h4f98,
// 16'h45a9, 16'h3a47, 16'h2dbf, 16'h2042,
// 16'h1226, 16'h03a5, 16'hf514, 16'he6bc,
// 16'hd8e5, 16'hcbdb, 16'hbfdf, 16'hb52f,
// 16'hac04, 16'ha48b, 16'h9ef1, 16'h9b46,
// 16'h99b1, 16'h9a21, 16'h9cb1, 16'ha137,
// 16'ha7b1, 16'haff0, 16'hb9d0, 16'hc51f,
// 16'hd19c, 16'hdf0a, 16'hed26, 16'hfb9d,
// 16'h0a34, 16'h188f, 16'h266d, 16'h3385,
// 16'h3f8e, 16'h4a52, 16'h538f, 16'h5b22,
// 16'h60d3, 16'h6496, 16'h664a, 16'h65ed,
// 16'h637f, 16'h5f0f, 16'h58ac, 16'h5086,
// 16'h46b4, 16'h3b7c, 16'h2f09, 16'h21a7,
// 16'h1393, 16'h051b, 16'hf687, 16'he827,
// 16'hda3e, 16'hcd20, 16'hc102, 16'hb632,
// 16'hacd9, 16'ha539, 16'h9f65, 16'h9b93,
// 16'h99bb, 16'h9a05, 16'h9c52, 16'ha0b0,
// 16'ha6f4, 16'haf09, 16'hb8c4, 16'hc3ee,
// 16'hd050, 16'hddaa, 16'hebb4, 16'hfa2d,
// 16'h08bd, 16'h1726, 16'h2510, 16'h3241,
// 16'h3e69, 16'h494d, 16'h52b9, 16'h5a70,
// 16'h605b, 16'h644c, 16'h6635, 16'h6610,
// 16'h63d4, 16'h5f95, 16'h596a, 16'h5164,
// 16'h47c6, 16'h3ca6, 16'h3056, 16'h2307,
// 16'h1520, 16'h0690, 16'hf7fc, 16'he990,
// 16'hdba0, 16'hce60, 16'hc22e, 16'hb733,
// 16'hadb8, 16'ha5e6, 16'h9fe6, 16'h9bdc,
// 16'h99d4, 16'h99e3, 16'h9c02, 16'ha028,
// 16'ha63e, 16'hae29, 16'hb7b7, 16'hc2c2,
// 16'hcf06, 16'hdc4c, 16'hea46, 16'hf8b9,
// 16'h0748, 16'h15b8, 16'h23b6, 16'h30f7,
// 16'h3d42, 16'h4844, 16'h51db, 16'h59c1,
// 16'h5fd7, 16'h6420, 16'h661a, 16'h662d,
// 16'h6425, 16'h6019, 16'h5a1c, 16'h5246,
// 16'h48cd, 16'h3dd3, 16'h319e, 16'h2463,
// 16'h1670, 16'h0801, 16'hf974, 16'heafb,
// 16'hdcfd, 16'hcfab, 16'hc355, 16'hb841,
// 16'hae93, 16'ha69e, 16'ha067, 16'h9c2c,
// 16'h99f2, 16'h99c8, 16'h9bb6, 16'h9fa5,
// 16'ha58e, 16'had49, 16'hb6b1, 16'hc199,
// 16'hcdbe, 16'hdaf0, 16'he8da, 16'hf742,
// 16'h05d6, 16'h1449, 16'h2257, 16'h2fb1,
// 16'h3c10, 16'h473f, 16'h50f5, 16'h590b,
// 16'h5f54, 16'h63a8, 16'h6601, 16'h6640,
// 16'h6471, 16'h6099, 16'h5ac8, 16'h5326,
// 16'h49ce, 16'h3eff, 16'h32df, 16'h25c4,
// 16'h17d6, 16'h097c, 16'hfae2, 16'hec70,
// 16'hde58, 16'hd0f5, 16'hc487, 16'hb949,
// 16'haf7d, 16'ha752, 16'ha0f2, 16'h9c80,
// 16'h9a14, 16'h99b5, 16'h9b6b, 16'h9f2c,
// 16'ha4df, 16'hac70, 16'hb5af, 16'hc071,
// 16'hcc7b, 16'hd994, 16'he76f, 16'hf5cf,
// 16'h0460, 16'h12db, 16'h20f7, 16'h2e61,
// 16'h3ae6, 16'h462c, 16'h5010, 16'h5852,
// 16'h5ec4, 16'h6357, 16'h65d6, 16'h6656,
// 16'h64b4, 16'h6114, 16'h5b73, 16'h53fc,
// 16'h4ad2, 16'h401f, 16'h3427, 16'h2719,
// 16'h1947, 16'h0ae9, 16'hfc5d, 16'hedd9,
// 16'hdfbe, 16'hd242, 16'hc5b7, 16'hba59,
// 16'hb067, 16'ha80d, 16'ha182, 16'h9cd9,
// 16'h9a3b, 16'h99a6, 16'h9b29, 16'h9eb3,
// 16'ha439, 16'hab98, 16'hb4b2, 16'hbf4d,
// 16'hcb3a, 16'hd83a, 16'he605, 16'hf45d,
// 16'h02e9, 16'h116d, 16'h1f92, 16'h2d17,
// 16'h39af, 16'h451c, 16'h4f24, 16'h5792,
// 16'h5e37, 16'h62f6, 16'h65b1, 16'h665e,
// 16'h64f8, 16'h6186, 16'h5c1a, 16'h54d0,
// 16'h4bcd, 16'h4145, 16'h3562, 16'h2875,
// 16'h1aad, 16'h0c5f, 16'hfdd1, 16'hef49,
// 16'he122, 16'hd390, 16'hc6ed, 16'hbb6c,
// 16'hb153, 16'ha8d1, 16'ha212, 16'h9d3b,
// 16'h9a65, 16'h999e, 16'h9ae9, 16'h9e44,
// 16'ha393, 16'haac9, 16'hb3b5, 16'hbe2e,
// 16'hc9fb, 16'hd6e4, 16'he49c, 16'hf2e9,
// 16'h0176, 16'h0ffa, 16'h1e30, 16'h2bc5,
// 16'h387a, 16'h4406, 16'h4e37, 16'h56cc,
// 16'h5da2, 16'h6295, 16'h6581, 16'h6667,
// 16'h6531, 16'h61f8, 16'h5cb7, 16'h55a4,
// 16'h4cc2, 16'h4265, 16'h369f, 16'h29cb,
// 16'h1c15, 16'h0dd1, 16'hff46, 16'hf0bc,
// 16'he284, 16'hd4e4, 16'hc822, 16'hbc87,
// 16'hb241, 16'ha999, 16'ha2a7, 16'h9da2,
// 16'h9a96, 16'h999a, 16'h9ab0, 16'h9dd7,
// 16'ha2f3, 16'ha9ff, 16'hb2bb, 16'hbd13,
// 16'hc8c0, 16'hd58c, 16'he337, 16'hf177,
// 16'hfffd, 16'h0e8e, 16'h1cc7, 16'h2a74,
// 16'h373f, 16'h42ef, 16'h4d42, 16'h5606,
// 16'h5d07, 16'h622d, 16'h654e, 16'h6667,
// 16'h656a, 16'h625d, 16'h5d5b, 16'h5665,
// 16'h4dbf, 16'h437b, 16'h37db, 16'h2b20,
// 16'h1d79, 16'h0f45, 16'h20b9, 16'hf231,
// 16'he3e8, 16'hd639, 16'hc95d, 16'hbd9e,
// 16'hb33b, 16'haa5f, 16'ha348, 16'h9e08,
// 16'h9acf, 16'h9999, 16'h9a7e, 16'h9d6d,
// 16'ha25e, 16'ha932, 16'hb1cc, 16'hbbf7,
// 16'hc788, 16'hd43a, 16'he1d1, 16'hf005,
// 16'hfe8b, 16'h0d17, 16'h1b63, 16'h291c,
// 16'h3606, 16'h41d1, 16'h4c4d, 16'h5534,
// 16'h5c6f, 16'h61ba, 16'h651a, 16'h6660,
// 16'h659c, 16'h62c3, 16'h5df0, 16'h572d,
// 16'h4eb0, 16'h4490, 16'h3918, 16'h2c69,
// 16'h1ee7, 16'h10ae, 16'h0235, 16'hf39f,
// 16'he552, 16'hd78e, 16'hca9b, 16'hbebc,
// 16'hb435, 16'hab2c, 16'ha3eb, 16'h9e76,
// 16'h9b0b, 16'h99a0, 16'h9a4f, 16'h9d0b,
// 16'ha1c9, 16'ha86e, 16'hb0dd, 16'hbae1,
// 16'hc652, 16'hd2ea, 16'he06d, 16'hee94,
// 16'hfd16, 16'h0ba4, 16'h19fa, 16'h27c7,
// 16'h34c4, 16'h40b5, 16'h4b4e, 16'h5467,
// 16'h5bc8, 16'h614b, 16'h64d9, 16'h6659,
// 16'h65c5, 16'h6328, 16'h5e7c, 16'h57f5,
// 16'h4f97, 16'h45a9, 16'h3a48, 16'h2dbd,
// 16'h2045, 16'h1223, 16'h03a7, 16'hf513,
// 16'he6bd, 16'hd8e3, 16'hcbde, 16'hbfdc,
// 16'hb530, 16'hac06, 16'ha488, 16'h9ef3,
// 16'h9b44, 16'h99b2, 16'h9a22, 16'h9cb1,
// 16'ha135, 16'ha7b3, 16'hafed, 16'hb9d5,
// 16'hc51b, 16'hd19d, 16'hdf0b, 16'hed23,
// 16'hfba1, 16'h0a32, 16'h188f, 16'h266e,
// 16'h3383, 16'h3f90, 16'h4a51, 16'h5391,
// 16'h5b20, 16'h60d4, 16'h6495, 16'h664b,
// 16'h65ed, 16'h6380, 16'h5f0d, 16'h58ae,
// 16'h5083, 16'h46b8, 16'h3b79, 16'h2f0b,
// 16'h21a6, 16'h1392, 16'h051d, 16'hf686,
// 16'he827, 16'hda40, 16'hcd1d, 16'hc104,
// 16'hb630, 16'hacdc, 16'ha536, 16'h9f69,
// 16'h9b8d, 16'h99c1, 16'h9a20, 16'h9c57,
// 16'ha0ab, 16'ha6f8, 16'haf07, 16'hb8c5,
// 16'hc3ed, 16'hd050, 16'hddaa, 16'hebb7,
// 16'hfa28, 16'h08c1, 16'h1722, 16'h2514,
// 16'h323e, 16'h3e6b, 16'h494c, 16'h52b9,
// 16'h5a71, 16'h605a, 16'h644c, 16'h6636,
// 16'h660f, 16'h63d5, 16'h5f96, 16'h5967,
// 16'h5167, 16'h47c3, 16'h3ca9, 16'h3056,
// 16'h2304, 16'h1503, 16'h068d, 16'hf7ff,
// 16'he990, 16'hdb9d, 16'hce63, 16'hc22b,
// 16'hb735, 16'hadb9, 16'ha5e4, 16'h9fe7,
// 16'h9bdb, 16'h99d4, 16'h99e6, 16'h9bfe,
// 16'ha02b, 16'ha63c, 16'hae2a, 16'hb7b7,
// 16'hc2c2, 16'hcf05, 16'hdc4d, 16'hea46,
// 16'hf8b8, 16'h0749, 16'h15b8, 16'h23b6,
// 16'h30f8, 16'h3d3f, 16'h4848, 16'h51d8,
// 16'h59c3, 16'h5fd6, 16'h6420, 16'h661b,
// 16'h662c, 16'h6425, 16'h601a, 16'h5a19,
// 16'h524b, 16'h48c8, 16'h3dd7, 16'h319b,
// 16'h2465, 16'h166d, 16'h0806, 16'hf96e,
// 16'heb20, 16'hdcfb, 16'hcfa9, 16'hc359,
// 16'hb83d, 16'hae97, 16'ha69b, 16'ha068,
// 16'h9c2d, 16'h99f0, 16'h99cc, 16'h9bb0,
// 16'h9fab, 16'ha58a, 16'had4b, 16'hb6b2,
// 16'hc196, 16'hcdc1, 16'hdaed, 16'he8dd,
// 16'hf740, 16'h05d7, 16'h144a, 16'h2254,
// 16'h2fb4, 16'h3c0d, 16'h4742, 16'h50f3,
// 16'h590c, 16'h5f53, 16'h63a9, 16'h6601,
// 16'h663f, 16'h6472, 16'h6098, 16'h5ac9,
// 16'h5326, 16'h49ce, 16'h3efe, 16'h32e1,
// 16'h25c1, 16'h17da, 16'h0978, 16'hfae5,
// 16'hec6d, 16'hde5a, 16'hd0f6, 16'hc484,
// 16'hb94c, 16'haf7a, 16'ha755, 16'ha0ef,
// 16'h9c84, 16'h9a0f, 16'h99ba, 16'h9b68,
// 16'h9f2c, 16'ha4e1, 16'hac6e, 16'hb5b1,
// 16'hc06f, 16'hcc7d, 16'hd992, 16'he771,
// 16'hf5ce, 16'h0460, 16'h12dc, 16'h20f4,
// 16'h2e65, 16'h3ae3, 16'h462d, 16'h5011,
// 16'h5850, 16'h5ec6, 16'h6354, 16'h65da,
// 16'h6652, 16'h64b9, 16'h6110, 16'h5b73,
// 16'h53fe, 16'h4acf, 16'h4023, 16'h3425,
// 16'h2718, 16'h1947, 16'h0aeb, 16'hfc5a,
// 16'heddc, 16'hdfbd, 16'hd240, 16'hc5ba,
// 16'hba58, 16'hb065, 16'ha811, 16'ha17e,
// 16'h9cdc, 16'h9a39, 16'h99a7, 16'h9b28,
// 16'h9eb5, 16'ha437, 16'hab9a, 16'hb4b0,
// 16'hbf4e, 16'hcb3a, 16'hd83b, 16'he604,
// 16'hf45e, 16'h02e7, 16'h1170, 16'h1f90,
// 16'h2d18, 16'h39ae, 16'h451d, 16'h4f24,
// 16'h5792, 16'h5e36, 16'h62f7, 16'h65b0,
// 16'h665f, 16'h64f7, 16'h6187, 16'h5c18,
// 16'h54d2, 16'h4bcc, 16'h4144, 16'h3565,
// 16'h2872, 16'h1aaf, 16'h0c5d, 16'hfdd2,
// 16'hef4a, 16'he120, 16'hd393, 16'hc6e9,
// 16'hbb6f, 16'hb153, 16'ha8ce, 16'ha215,
// 16'h9d3a, 16'h9a65, 16'h999f, 16'h9ae8,
// 16'h9e43, 16'ha395, 16'haac8, 16'hb3b6,
// 16'hbe2b, 16'hca20, 16'hd6de, 16'he4a1,
// 16'hf2e6, 16'h0176, 16'h0ffc, 16'h1e2e,
// 16'h2bc6, 16'h3878, 16'h4409, 16'h4e34,
// 16'h56cf, 16'h5da0, 16'h6295, 16'h6581,
// 16'h6668, 16'h6531, 16'h61f6, 16'h5cba,
// 16'h559f, 16'h4cc8, 16'h4260, 16'h36a3,
// 16'h29c8, 16'h1c15, 16'h0dd3, 16'hff43,
// 16'hf0c0, 16'he282, 16'hd4e3, 16'hc825,
// 16'hbc82, 16'hb247, 16'ha994, 16'ha2aa,
// 16'h9da1, 16'h9a95, 16'h999c, 16'h9aaf,
// 16'h9dd5, 16'ha2f8, 16'ha9f9, 16'hb2c0,
// 16'hbd10, 16'hc8c1, 16'hd58d, 16'he336,
// 16'hf176, 16'h2020, 16'h0e8b, 16'h1cc9,
// 16'h2a72, 16'h3740, 16'h42ef, 16'h4d43,
// 16'h5603, 16'h5d0c, 16'h6227, 16'h6553,
// 16'h6664, 16'h656b, 16'h625f, 16'h5d57,
// 16'h5669, 16'h4dbd, 16'h437a, 16'h37e0,
// 16'h2b18, 16'h1d81, 16'h0f3f, 16'h20bd,
// 16'hf22e, 16'he3ea, 16'hd638, 16'hc95e,
// 16'hbd9e, 16'hb33a, 16'haa60, 16'ha346,
// 16'h9e0b, 16'h9acd, 16'h999a, 16'h9a7e,
// 16'h9d6d, 16'ha25c, 16'ha936, 16'hb1c6,
// 16'hbbfd, 16'hc784, 16'hd43d, 16'he1cf,
// 16'hf006, 16'hfe88, 16'h0d1b, 16'h1b60,
// 16'h2920, 16'h3601, 16'h41d6, 16'h4c47,
// 16'h553b, 16'h5c69, 16'h61bf, 16'h6516,
// 16'h6662, 16'h659b, 16'h62c5, 16'h5ded,
// 16'h5731, 16'h4eab, 16'h4495, 16'h3912,
// 16'h2c71, 16'h1edf, 16'h10b4, 16'h0231,
// 16'hf39f, 16'he555, 16'hd78c, 16'hca9b,
// 16'hbebd, 16'hb432, 16'hab30, 16'ha3e7,
// 16'h9e7a, 16'h9b08, 16'h99a2, 16'h9a4e,
// 16'h9d0b, 16'ha1c9, 16'ha86f, 16'hb0db,
// 16'hbae4, 16'hc650, 16'hd2eb, 16'he06d,
// 16'hee93, 16'hfd16, 16'h0ba5, 16'h19fa,
// 16'h27c6, 16'h34c5, 16'h40b4, 16'h4b4d,
// 16'h546b, 16'h5bc3, 16'h6150, 16'h64d5,
// 16'h665b, 16'h65c6, 16'h6325, 16'h5e80,
// 16'h57f1, 16'h4f9b, 16'h45a6, 16'h3a49,
// 16'h2dbe, 16'h2043, 16'h1225, 16'h03a6,
// 16'hf513, 16'he6bd, 16'hd8e3, 16'hcbdf,
// 16'hbfda, 16'hb534, 16'hac20, 16'ha48e,
// 16'h9eee, 16'h9b49, 16'h99ae, 16'h9a25,
// 16'h9cad, 16'ha13a, 16'ha7ad, 16'haff4,
// 16'hb9cf, 16'hc51f, 16'hd19b, 16'hdf0b,
// 16'hed24, 16'hfba0, 16'h0a33, 16'h188f,
// 16'h266d, 16'h3385, 16'h3f8d, 16'h4a53,
// 16'h5391, 16'h5b1e, 16'h60d7, 16'h6493,
// 16'h664c, 16'h65ec, 16'h6380, 16'h5f0d,
// 16'h58ae, 16'h5085, 16'h46b4, 16'h3b7d,
// 16'h2f08, 16'h21a7, 16'h1393, 16'h051a,
// 16'hf689, 16'he826, 16'hda3e, 16'hcd21,
// 16'hc120, 16'hb633, 16'hacdb, 16'ha535,
// 16'h9f6a, 16'h9b8e, 16'h99bf, 16'h9a02,
// 16'h9c54, 16'ha0af, 16'ha6f4, 16'haf0a,
// 16'hb8c4, 16'hc3ec, 16'hd052, 16'hdda9,
// 16'hebb5, 16'hfa2d, 16'h08bc, 16'h1726,
// 16'h2512, 16'h323e, 16'h3e6b, 16'h494d,
// 16'h52b8, 16'h5a72, 16'h6059, 16'h644c,
// 16'h6637, 16'h660f, 16'h63d3, 16'h5f99,
// 16'h5963, 16'h516c, 16'h47bf, 16'h3cab,
// 16'h3054, 16'h2307, 16'h14ff, 16'h0692,
// 16'hf7f9, 16'he995, 16'hdb9a, 16'hce65,
// 16'hc229, 16'hb738, 16'hadb5, 16'ha5e8,
// 16'h9fe5, 16'h9bda, 16'h99d8, 16'h99df,
// 16'h9c07, 16'ha022, 16'ha644, 16'hae24,
// 16'hb7ba, 16'hc2c1, 16'hcf06, 16'hdc4b,
// 16'hea49, 16'hf8b5, 16'h074b, 16'h15b7,
// 16'h23b6, 16'h30f8, 16'h3d40, 16'h4847,
// 16'h51d9, 16'h59c1, 16'h5fd8, 16'h63ff,
// 16'h661c, 16'h662c, 16'h6424, 16'h601b,
// 16'h5a18, 16'h524c, 16'h48c7, 16'h3dd9,
// 16'h3199, 16'h2467, 16'h166b, 16'h0807,
// 16'hf96f, 16'heaff, 16'hdcfb, 16'hcfaa,
// 16'hc357, 16'hb83f, 16'hae96, 16'ha69b,
// 16'ha069, 16'h9c2c, 16'h99f0, 16'h99cb,
// 16'h9bb3, 16'h9fa7, 16'ha58f, 16'had46,
// 16'hb6b5, 16'hc194, 16'hcdc2, 16'hdaee,
// 16'he8db, 16'hf742, 16'h05d5, 16'h144b,
// 16'h2254, 16'h2fb3, 16'h3c0f, 16'h473f,
// 16'h50f6, 16'h590a, 16'h5f53, 16'h63ab,
// 16'h65fe, 16'h6642, 16'h6470, 16'h6099,
// 16'h5ac8, 16'h5326, 16'h49d0, 16'h3efb,
// 16'h32e4, 16'h25be, 16'h17dc, 16'h0977,
// 16'hfae6, 16'hec6d, 16'hde5a, 16'hd0f5,
// 16'hc487, 16'hb947, 16'haf80, 16'ha750,
// 16'ha0f3, 16'h9c80, 16'h9a14, 16'h99b4,
// 16'h9b6d, 16'h9f2a, 16'ha4df, 16'hac72,
// 16'hb5ad, 16'hc071, 16'hcc7d, 16'hd990,
// 16'he774, 16'hf5cb, 16'h0462, 16'h12db,
// 16'h20f5, 16'h2e65, 16'h3ae2, 16'h462e,
// 16'h5011, 16'h584e, 16'h5eca, 16'h6350,
// 16'h65dd, 16'h6650, 16'h64b9, 16'h6110,
// 16'h5b74, 16'h53fd, 16'h4ad1, 16'h4020,
// 16'h3427, 16'h2718, 16'h1947, 16'h0aea,
// 16'hfc5c, 16'hedda, 16'hdfbd, 16'hd243,
// 16'hc5b6, 16'hba5a, 16'hb066, 16'ha80d,
// 16'ha183, 16'h9cd9, 16'h9a3a, 16'h99a7,
// 16'h9b28, 16'h9eb4, 16'ha438, 16'hab9a,
// 16'hb4af, 16'hbf4f, 16'hcb3a, 16'hd839,
// 16'he607, 16'hf45a, 16'h02ec, 16'h116b,
// 16'h1f95, 16'h2d13, 16'h39b2, 16'h451b,
// 16'h4f25, 16'h5791, 16'h5e38, 16'h62f4,
// 16'h65b3, 16'h665d, 16'h64f8, 16'h6187,
// 16'h5c18, 16'h54d1, 16'h4bcd, 16'h4143,
// 16'h3566, 16'h2871, 16'h1aaf, 16'h0c5e,
// 16'hfdd1, 16'hef4a, 16'he122, 16'hd38e,
// 16'hc6f0, 16'hbb69, 16'hb156, 16'ha8ce,
// 16'ha214, 16'h9d3b, 16'h9a64, 16'h999f,
// 16'h9ae8, 16'h9e45, 16'ha392, 16'haacb,
// 16'hb3b3, 16'hbe2f, 16'hc9fa, 16'hd6e5,
// 16'he49b, 16'hf2eb, 16'h0174, 16'h0ffb,
// 16'h1e2f, 16'h2bc6, 16'h3879, 16'h4407,
// 16'h4e37, 16'h56cb, 16'h5da3, 16'h6295,
// 16'h657f, 16'h666a, 16'h652f, 16'h61f8,
// 16'h5cb9, 16'h55a0, 16'h4cc6, 16'h4262,
// 16'h36a1, 16'h29cb, 16'h1c13, 16'h0dd4,
// 16'hff42, 16'hf0c0, 16'he281, 16'hd4e7,
// 16'hc820, 16'hbc87, 16'hb241, 16'ha999,
// 16'ha2a7, 16'h9da3, 16'h9a94, 16'h999b,
// 16'h9ab0, 16'h9dd6, 16'ha2f5, 16'ha9fd,
// 16'hb2bd, 16'hbd12, 16'hc8bf, 16'hd58e,
// 16'he336, 16'hf178, 16'hfffe, 16'h0e8c,
// 16'h1cc7, 16'h2a74, 16'h3740, 16'h42ee,
// 16'h4d44, 16'h5603, 16'h5d09, 16'h622d,
// 16'h654c, 16'h666a, 16'h6567, 16'h6261,
// 16'h5d56, 16'h566a, 16'h4dbb, 16'h437c,
// 16'h37de, 16'h2b1a, 16'h1d7f, 16'h0f41,
// 16'h20bb, 16'hf230, 16'he3e8, 16'hd63a,
// 16'hc95c, 16'hbda0, 16'hb339, 16'haa60,
// 16'ha346, 16'h9e0b, 16'h9acd, 16'h999b,
// 16'h9a7c, 16'h9d6f, 16'ha25a, 16'ha937,
// 16'hb1c7, 16'hbbfb, 16'hc786, 16'hd43a,
// 16'he1d2, 16'hf004, 16'hfe8a, 16'h0d1a,
// 16'h1b5f, 16'h2921, 16'h3601, 16'h41d4,
// 16'h4c4b, 16'h5537, 16'h5c6c, 16'h61bc,
// 16'h6519, 16'h665f, 16'h659f, 16'h62c1,
// 16'h5df0, 16'h572f, 16'h4ead, 16'h4494,
// 16'h3913, 16'h2c6f, 16'h1ee0, 16'h10b5,
// 16'h0230, 16'hf3a1, 16'he551, 16'hd78f,
// 16'hca99, 16'hbec0, 16'hb42f, 16'hab33,
// 16'ha3e4, 16'h9e7b, 16'h9b08, 16'h99a2,
// 16'h9a4e, 16'h9d0c, 16'ha1c7, 16'ha870,
// 16'hb0db, 16'hbae4, 16'hc64f, 16'hd2ed,
// 16'he06a, 16'hee96, 16'hfd15, 16'h0ba4,
// 16'h19fb, 16'h27c5, 16'h34c7, 16'h40b2,
// 16'h4b4f, 16'h5468, 16'h5bc6, 16'h614e,
// 16'h64d6, 16'h665b, 16'h65c5, 16'h6326,
// 16'h5e7f, 16'h57f1, 16'h4f9d, 16'h45a3,
// 16'h3a4c, 16'h2dba, 16'h2048, 16'h1221,
// 16'h03a9, 16'hf510, 16'he6bf, 16'hd8e3,
// 16'hcbdd, 16'hbfde, 16'hb52f, 16'hac04,
// 16'ha48b, 16'h9ef0, 16'h9b48, 16'h99ae,
// 16'h9a26, 16'h9cac, 16'ha13a, 16'ha7af,
// 16'haff0, 16'hb9d3, 16'hc51c, 16'hd19e,
// 16'hdf08, 16'hed27, 16'hfb9e, 16'h0a33,
// 16'h188f, 16'h266e, 16'h3383, 16'h3f91,
// 16'h4a4e, 16'h5394, 16'h5b1d, 16'h60d7,
// 16'h6494, 16'h664a, 16'h65ee, 16'h637f,
// 16'h5f0d, 16'h58af, 16'h5084, 16'h46b4,
// 16'h3b7e, 16'h2f05, 16'h21ab, 16'h1390,
// 16'h051d, 16'hf686, 16'he827, 16'hda3f,
// 16'hcd1f, 16'hc102, 16'hb632, 16'hacda,
// 16'ha537, 16'h9f69, 16'h9b8c, 16'h99c3,
// 16'h99fe, 16'h9c57, 16'ha0ae, 16'ha6f3,
// 16'haf0c, 16'hb8c1, 16'hc3f0, 16'hd04e,
// 16'hddad, 16'hebb3, 16'hfa2c, 16'h08be,
// 16'h1724, 16'h2513, 16'h3240, 16'h3e68,
// 16'h494f, 16'h52b5, 16'h5a76, 16'h6055,
// 16'h6451, 16'h6631, 16'h6613, 16'h63d2,
// 16'h5f98, 16'h5965, 16'h5169, 16'h47c2,
// 16'h3caa, 16'h3054, 16'h2305, 16'h1504,
// 16'h068c, 16'hf820, 16'he98d, 16'hdba0,
// 16'hce62, 16'hc22b, 16'hb736, 16'hadb6,
// 16'ha5e7, 16'h9fe7, 16'h9bd8, 16'h99d8,
// 16'h99e2, 16'h9c02, 16'ha028, 16'ha63e,
// 16'hae27, 16'hb7bb, 16'hc2be, 16'hcf09,
// 16'hdc49, 16'hea49, 16'hf8b6, 16'h074a,
// 16'h15b7, 16'h23b7, 16'h30f6, 16'h3d42,
// 16'h4846, 16'h51d8, 16'h59c4, 16'h5fd4,
// 16'h6403, 16'h6618, 16'h662e, 16'h6424,
// 16'h6019, 16'h5a1d, 16'h5245, 16'h48cd,
// 16'h3dd4, 16'h319c, 16'h2466, 16'h166c,
// 16'h0806, 16'hf96f, 16'heaff, 16'hdcfb,
// 16'hcfaa, 16'hc358, 16'hb83d, 16'hae98,
// 16'ha699, 16'ha06a, 16'h9c2b, 16'h99f2,
// 16'h99c9, 16'h9bb5, 16'h9fa6, 16'ha58e,
// 16'had48, 16'hb6b3, 16'hc197, 16'hcdc0,
// 16'hdaef, 16'he8d9, 16'hf744, 16'h05d5,
// 16'h1449, 16'h2258, 16'h2fae, 16'h3c13,
// 16'h473d, 16'h50f6, 16'h590b, 16'h5f53,
// 16'h63a9, 16'h6602, 16'h663d, 16'h6474,
// 16'h6097, 16'h5ac8, 16'h5329, 16'h49ca,
// 16'h3f01, 16'h32e0, 16'h25c0, 16'h17dc,
// 16'h0975, 16'hfae9, 16'hec69, 16'hde5d,
// 16'hd0f4, 16'hc487, 16'hb948, 16'haf7e,
// 16'ha752, 16'ha0f1, 16'h9c83, 16'h9a10,
// 16'h99b8, 16'h9b6a, 16'h9f2c, 16'ha4df,
// 16'hac70, 16'hb5af, 16'hc070, 16'hcc7d,
// 16'hd992, 16'he770, 16'hf5cf, 16'h045f,
// 16'h12dd, 16'h20f4, 16'h2e65, 16'h3ae1,
// 16'h4631, 16'h500d, 16'h5852, 16'h5ec6,
// 16'h6354, 16'h65d9, 16'h6655, 16'h64b3,
// 16'h6116, 16'h5b70, 16'h53ff, 16'h4acf,
// 16'h4023, 16'h3424, 16'h271b, 16'h1944,
// 16'h0aeb, 16'hfc5d, 16'hedda, 16'hdfbd,
// 16'hd242, 16'hc5b6, 16'hba5c, 16'hb064,
// 16'ha810, 16'ha17f, 16'h9cdb, 16'h9a3b,
// 16'h99a5, 16'h9b2a, 16'h9eb1, 16'ha43c,
// 16'hab96, 16'hb4b3, 16'hbf4b, 16'hcb3c,
// 16'hd839, 16'he607, 16'hf45a, 16'h02eb,
// 16'h116d, 16'h1f91, 16'h2d18, 16'h39ae,
// 16'h451d, 16'h4f25, 16'h5790, 16'h5e38,
// 16'h62f5, 16'h65b2, 16'h665e, 16'h64f8,
// 16'h6185, 16'h5c1a, 16'h54d0, 16'h4bce,
// 16'h4143, 16'h3564, 16'h2874, 16'h1aac,
// 16'h0c61, 16'hfdce, 16'hef4d, 16'he11f,
// 16'hd392, 16'hc6eb, 16'hbb6f, 16'hb150,
// 16'ha8d3, 16'ha210, 16'h9d3d, 16'h9a65,
// 16'h999d, 16'h9aea, 16'h9e41, 16'ha397,
// 16'haac7, 16'hb3b5, 16'hbe2f, 16'hc9f9,
// 16'hd6e6, 16'he49b, 16'hf2e9, 16'h0175,
// 16'h0ffc, 16'h1e2f, 16'h2bc5, 16'h3879,
// 16'h4407, 16'h4e37, 16'h56cb, 16'h5da5,
// 16'h6290, 16'h6585, 16'h6664, 16'h6533,
// 16'h61f7, 16'h5cb8, 16'h55a1, 16'h4cc6,
// 16'h4261, 16'h36a2, 16'h29cb, 16'h1c12,
// 16'h0dd5, 16'hff42, 16'hf0bf, 16'he284,
// 16'hd4e3, 16'hc824, 16'hbc83, 16'hb245,
// 16'ha996, 16'ha2aa, 16'h9da0, 16'h9a97,
// 16'h9999, 16'h9ab1, 16'h9dd5, 16'ha2f6,
// 16'ha9fd, 16'hb2bc, 16'hbd13, 16'hc8bf,
// 16'hd58d, 16'he337, 16'hf176, 16'h2020,
// 16'h0e8b, 16'h1cc8, 16'h2a73, 16'h3740,
// 16'h42ef, 16'h4d42, 16'h5605, 16'h5d09,
// 16'h622a, 16'h6551, 16'h6665, 16'h656a,
// 16'h6260, 16'h5d56, 16'h566a, 16'h4dbc,
// 16'h437b, 16'h37de, 16'h2b1b, 16'h1d7e,
// 16'h0f41, 16'h20bc, 16'hf22f, 16'he3e9,
// 16'hd638, 16'hc95e, 16'hbd9f, 16'hb33a,
// 16'haa5f, 16'ha347, 16'h9e0a, 16'h9acd,
// 16'h999c, 16'h9a7a, 16'h9d71, 16'ha25b,
// 16'ha933, 16'hb1cc, 16'hbbf7, 16'hc787,
// 16'hd43d, 16'he1cd, 16'hf009, 16'hfe87,
// 16'h0d1a, 16'h1b62, 16'h291c, 16'h3607,
// 16'h41cf, 16'h4c4e, 16'h5536, 16'h5c6a,
// 16'h61c1, 16'h6513, 16'h6665, 16'h6599,
// 16'h62c6, 16'h5dec, 16'h5732, 16'h4eac,
// 16'h4492, 16'h3917, 16'h2c6b, 16'h1ee4,
// 16'h10b2, 16'h0231, 16'hf3a1, 16'he552,
// 16'hd78e, 16'hca9a, 16'hbebe, 16'hb432,
// 16'hab2f, 16'ha3e8, 16'h9e79, 16'h9b08,
// 16'h99a3, 16'h9a4c, 16'h9d0e, 16'ha1c5,
// 16'ha872, 16'hb0d9, 16'hbae5, 16'hc64f,
// 16'hd2ed, 16'he069, 16'hee98, 16'hfd12,
// 16'h0ba7, 16'h19f9, 16'h27c6, 16'h34c7,
// 16'h40b1, 16'h4b51, 16'h5466, 16'h5bc7,
// 16'h614d, 16'h64d7, 16'h665b, 16'h65c4,
// 16'h6328, 16'h5e7c, 16'h57f5, 16'h4f98,
// 16'h45a7, 16'h3a49, 16'h2dbe, 16'h2042,
// 16'h1228, 16'h03a1, 16'hf518, 16'he6b9,
// 16'hd8e7, 16'hcbda, 16'hbfdf, 16'hb530,
// 16'hac02, 16'ha48e, 16'h9eed, 16'h9b49,
// 16'h99af, 16'h9a24, 16'h9cae, 16'ha138,
// 16'ha7b0, 16'haff1, 16'hb9d1, 16'hc51e,
// 16'hd19b, 16'hdf0c, 16'hed23, 16'hfba1,
// 16'h0a31, 16'h1891, 16'h266c, 16'h3385,
// 16'h3f8e, 16'h4a52, 16'h5391, 16'h5b1f,
// 16'h60d5, 16'h6495, 16'h664a, 16'h65ee,
// 16'h637e, 16'h5f0f, 16'h58ad, 16'h5085,
// 16'h46b4, 16'h3b7d, 16'h2f08, 16'h21a7,
// 16'h1394, 16'h0518, 16'hf68c, 16'he821,
// 16'hda44, 16'hcd1b, 16'hc105, 16'hb630,
// 16'hacdb, 16'ha536, 16'h9f69, 16'h9b8f,
// 16'h99bf, 16'h9a02, 16'h9c53, 16'ha0b1,
// 16'ha6f1, 16'haf0f, 16'hb8be, 16'hc3f2,
// 16'hd04d, 16'hddac, 16'hebb4, 16'hfa2d,
// 16'h08bb, 16'h1728, 16'h250f, 16'h3242,
// 16'h3e67, 16'h494f, 16'h52b6, 16'h5a75,
// 16'h6056, 16'h644f, 16'h6634, 16'h6610,
// 16'h63d5, 16'h5f95, 16'h5968, 16'h5167,
// 16'h47c3, 16'h3ca9, 16'h3055, 16'h2305,
// 16'h1503, 16'h068c, 16'hf820, 16'he98f,
// 16'hdb9d, 16'hce64, 16'hc229, 16'hb738,
// 16'hadb6, 16'ha5e6, 16'h9fe7, 16'h9bd9,
// 16'h99d8, 16'h99e0, 16'h9c05, 16'ha025,
// 16'ha641, 16'hae26, 16'hb7b9, 16'hc2c1,
// 16'hcf06, 16'hdc4c, 16'hea48, 16'hf8b6,
// 16'h0749, 16'h15b9, 16'h23b4, 16'h30fb,
// 16'h3d3d, 16'h484a, 16'h51d5, 16'h59c6,
// 16'h5fd3, 16'h6403, 16'h661a, 16'h662b,
// 16'h6426, 16'h6019, 16'h5a1b, 16'h5249,
// 16'h48c9, 16'h3dd6, 16'h319c, 16'h2464,
// 16'h166f, 16'h0802, 16'hf973, 16'heafc,
// 16'hdcfd, 16'hcfa9, 16'hc358, 16'hb83e,
// 16'hae96, 16'ha69b, 16'ha06a, 16'h9c2a,
// 16'h99f4, 16'h99c6, 16'h9bb7, 16'h9fa5,
// 16'ha58e, 16'had49, 16'hb6b2, 16'hc197,
// 16'hcdc0, 16'hdaee, 16'he8db, 16'hf744,
// 16'h05d3, 16'h144b, 16'h2257, 16'h2fae,
// 16'h3c15, 16'h473b, 16'h50f6, 16'h590d,
// 16'h5f50, 16'h63ac, 16'h65ff, 16'h6640,
// 16'h6473, 16'h6095, 16'h5acc, 16'h5323,
// 16'h49d0, 16'h3eff, 16'h32de, 16'h25c4,
// 16'h17d7, 16'h097a, 16'hfae5, 16'hec6c,
// 16'hde5b, 16'hd0f5, 16'hc486, 16'hb94a,
// 16'haf7b, 16'ha755, 16'ha0ef, 16'h9c84,
// 16'h9a0f, 16'h99b9, 16'h9b69, 16'h9f2d,
// 16'ha4df, 16'hac70, 16'hb5ae, 16'hc071,
// 16'hcc7c, 16'hd993, 16'he771, 16'hf5cd,
// 16'h0461, 16'h12da, 16'h20f7, 16'h2e63,
// 16'h3ae4, 16'h462d, 16'h5011, 16'h584e,
// 16'h5eca, 16'h6351, 16'h65db, 16'h6653,
// 16'h64b6, 16'h6113, 16'h5b73, 16'h53fc,
// 16'h4ad1, 16'h4022, 16'h3424, 16'h271c,
// 16'h1942, 16'h0aee, 16'hfc59, 16'heddd,
// 16'hdfbb, 16'hd243, 16'hc5b7, 16'hba5a,
// 16'hb064, 16'ha811, 16'ha17e, 16'h9cdd,
// 16'h9a39, 16'h99a5, 16'h9b2a, 16'h9eb2,
// 16'ha43b, 16'hab96, 16'hb4b4, 16'hbf49,
// 16'hcb3f, 16'hd835, 16'he60b, 16'hf456,
// 16'h02f0, 16'h1167, 16'h1f98, 16'h2d11,
// 16'h39b3, 16'h451b, 16'h4f25, 16'h5792,
// 16'h5e35, 16'h62f8, 16'h65b0, 16'h665f,
// 16'h64f8, 16'h6185, 16'h5c1a, 16'h54d0,
// 16'h4bce, 16'h4143, 16'h3566, 16'h2870,
// 16'h1ab0, 16'h0c5d, 16'hfdd2, 16'hef4b,
// 16'he120, 16'hd38f, 16'hc6ef, 16'hbb6b,
// 16'hb154, 16'ha8d1, 16'ha210, 16'h9d3e,
// 16'h9a63, 16'h999f, 16'h9ae9, 16'h9e42,
// 16'ha395, 16'haac9, 16'hb3b3, 16'hbe31,
// 16'hc9f8, 16'hd6e5, 16'he49c, 16'hf2e9,
// 16'h0175, 16'h0ffd, 16'h1e2d, 16'h2bc6,
// 16'h3879, 16'h4408, 16'h4e35, 16'h56ce,
// 16'h5da1, 16'h6294, 16'h6583, 16'h6664,
// 16'h6536, 16'h61f2, 16'h5cbd, 16'h559d,
// 16'h4cc9, 16'h425f, 16'h36a5, 16'h29c6,
// 16'h1c17, 16'h0dd1, 16'hff45, 16'hf0bd,
// 16'he284, 16'hd4e3, 16'hc825, 16'hbc81,
// 16'hb247, 16'ha994, 16'ha2ab, 16'h9da0,
// 16'h9a96, 16'h999a, 16'h9ab0, 16'h9dd6,
// 16'ha2f6, 16'ha9fc, 16'hb2bd, 16'hbd11,
// 16'hc8c2, 16'hd58b, 16'he339, 16'hf174,
// 16'h2020, 16'h0e8c, 16'h1cc8, 16'h2a73,
// 16'h3740, 16'h42ee, 16'h4d43, 16'h5605,
// 16'h5d08, 16'h622c, 16'h654e, 16'h6667,
// 16'h656a, 16'h625f, 16'h5d56, 16'h566b,
// 16'h4dba, 16'h437e, 16'h37db, 16'h2b1d,
// 16'h1d7d, 16'h0f41, 16'h20be, 16'hf22b,
// 16'he3ed, 16'hd636, 16'hc95e, 16'hbd9f,
// 16'hb339, 16'haa61, 16'ha346, 16'h9e0a,
// 16'h9acd, 16'h999b, 16'h9a7d, 16'h9d6e,
// 16'ha25b, 16'ha936, 16'hb1c8, 16'hbbfa,
// 16'hc787, 16'hd439, 16'he1d3, 16'hf003,
// 16'hfe8b, 16'h0d19, 16'h1b60, 16'h2921,
// 16'h3620, 16'h41d6, 16'h4c49, 16'h5538,
// 16'h5c6b, 16'h61be, 16'h6516, 16'h6663,
// 16'h659a, 16'h62c5, 16'h5dee, 16'h572f,
// 16'h4eae, 16'h4492, 16'h3915, 16'h2c6e,
// 16'h1ee1, 16'h10b3, 16'h0232, 16'hf3a0,
// 16'he552, 16'hd78e, 16'hca9a, 16'hbebf,
// 16'hb430, 16'hab32, 16'ha3e4, 16'h9e7d,
// 16'h9b07, 16'h99a1, 16'h9a50, 16'h9d08,
// 16'ha1cc, 16'ha86c, 16'hb0de, 16'hbae1,
// 16'hc653, 16'hd2e8, 16'he06e, 16'hee94,
// 16'hfd15, 16'h0ba5, 16'h19fa, 16'h27c7,
// 16'h34c4, 16'h40b4, 16'h4b4f, 16'h5466,
// 16'h5bc9, 16'h614b, 16'h64d9, 16'h6659,
// 16'h65c6, 16'h6325, 16'h5e80, 16'h57f2,
// 16'h4f99, 16'h45a8, 16'h3a48, 16'h2dbd,
// 16'h2046, 16'h1221, 16'h03a9, 16'hf511,
// 16'he6be, 16'hd8e4, 16'hcbdd, 16'hbfdd,
// 16'hb530, 16'hac02, 16'ha48f, 16'h9eec,
// 16'h9b4b, 16'h99ac, 16'h9a26, 16'h9cae,
// 16'ha137, 16'ha7b1, 16'haff0, 16'hb9d1,
// 16'hc520, 16'hd199, 16'hdf0c, 16'hed24,
// 16'hfba0, 16'h0a33, 16'h188e, 16'h266e,
// 16'h3384, 16'h3f90, 16'h4a50, 16'h5392,
// 16'h5b1e, 16'h60d6, 16'h6495, 16'h664a,
// 16'h65ee, 16'h637e, 16'h5f0e, 16'h58af,
// 16'h5083, 16'h46b6, 16'h3b7b, 16'h2f09,
// 16'h21a8, 16'h1391, 16'h051d, 16'hf685,
// 16'he829, 16'hda3d, 16'hcd20, 16'hc101,
// 16'hb633, 16'hacda, 16'ha536, 16'h9f69,
// 16'h9b8e, 16'h99bf, 16'h9a04, 16'h9c51,
// 16'ha0b2, 16'ha6f0, 16'haf0e, 16'hb8c0,
// 16'hc3f1, 16'hd04d, 16'hddad, 16'hebb2,
// 16'hfa2d, 16'h08bf, 16'h1723, 16'h2513,
// 16'h323f, 16'h3e68, 16'h4951, 16'h52b5,
// 16'h5a73, 16'h6059, 16'h644c, 16'h6637,
// 16'h660e, 16'h63d5, 16'h5f96, 16'h5967,
// 16'h5168, 16'h47c2, 16'h3caa, 16'h3054,
// 16'h2306, 16'h1502, 16'h068f, 16'hf7fc,
// 16'he992, 16'hdb9c, 16'hce63, 16'hc22c,
// 16'hb734, 16'hadb9, 16'ha5e5, 16'h9fe6,
// 16'h9bdb, 16'h99d4, 16'h99e6, 16'h9bff,
// 16'ha02a, 16'ha63c, 16'hae2a, 16'hb7b7,
// 16'hc2c3, 16'hcf04, 16'hdc4d, 16'hea46,
// 16'hf8b9, 16'h0747, 16'h15bb, 16'h23b2,
// 16'h30fb, 16'h3d3f, 16'h4846, 16'h51da,
// 16'h59c2, 16'h5fd6, 16'h6420, 16'h661c,
// 16'h662a, 16'h6427, 16'h6018, 16'h5a1b,
// 16'h5249, 16'h48ca, 16'h3dd5, 16'h319c,
// 16'h2465, 16'h166d, 16'h0806, 16'hf96e,
// 16'heb01, 16'hdcf8, 16'hcfad, 16'hc356,
// 16'hb83d, 16'hae9a, 16'ha696, 16'ha06d,
// 16'h9c2a, 16'h99f0, 16'h99cc, 16'h9bb2,
// 16'h9fa8, 16'ha58d, 16'had49, 16'hb6b2,
// 16'hc197, 16'hcdc1, 16'hdaed, 16'he8dc,
// 16'hf742, 16'h05d5, 16'h144a, 16'h2257,
// 16'h2fae, 16'h3c14, 16'h473c, 16'h50f6,
// 16'h590b, 16'h5f53, 16'h63aa, 16'h65ff,
// 16'h6641, 16'h6470, 16'h609a, 16'h5ac7,
// 16'h5326, 16'h49d0, 16'h3efc, 16'h32e3,
// 16'h25bf, 16'h17db, 16'h0978, 16'hfae5,
// 16'hec6d, 16'hde5a, 16'hd0f6, 16'hc486,
// 16'hb949, 16'haf7d, 16'ha751, 16'ha0f3,
// 16'h9c81, 16'h9a13, 16'h99b4, 16'h9b6d,
// 16'h9f29, 16'ha4e3, 16'hac6d, 16'hb5b0,
// 16'hc070, 16'hcc7d, 16'hd991, 16'he772,
// 16'hf5ce, 16'h045f, 16'h12dd, 16'h20f3,
// 16'h2e67, 16'h3ae0, 16'h4631, 16'h500d,
// 16'h5851, 16'h5ec9, 16'h6350, 16'h65dd,
// 16'h6651, 16'h64b8, 16'h6110, 16'h5b76,
// 16'h53fa, 16'h4ad3, 16'h4020, 16'h3426,
// 16'h2719, 16'h1946, 16'h0aea, 16'hfc5c,
// 16'heddc, 16'hdfbb, 16'hd244, 16'hc5b5,
// 16'hba5b, 16'hb066, 16'ha80d, 16'ha183,
// 16'h9cd8, 16'h9a3c, 16'h99a6, 16'h9b27,
// 16'h9eb5, 16'ha438, 16'hab9a, 16'hb4af,
// 16'hbf4f, 16'hcb39, 16'hd83b, 16'he605,
// 16'hf45c, 16'h02e9, 16'h116e, 16'h1f92,
// 16'h2d16, 16'h39af, 16'h451e, 16'h4f22,
// 16'h5794, 16'h5e35, 16'h62f7, 16'h65b0,
// 16'h6660, 16'h64f6, 16'h6188, 16'h5c17,
// 16'h54d2, 16'h4bcc, 16'h4144, 16'h3565,
// 16'h2872, 16'h1aae, 16'h0c60, 16'hfdcd,
// 16'hef4f, 16'he11c, 16'hd395, 16'hc6e9,
// 16'hbb70, 16'hb150, 16'ha8d2, 16'ha212,
// 16'h9d3b, 16'h9a66, 16'h999c, 16'h9aec,
// 16'h9e40, 16'ha396, 16'haac9, 16'hb3b3,
// 16'hbe30, 16'hc9f9, 16'hd6e6, 16'he49a,
// 16'hf2ec, 16'h0172, 16'h0ffe, 16'h1e2d,
// 16'h2bc7, 16'h3878, 16'h4408, 16'h4e36,
// 16'h56cb, 16'h5da6, 16'h628f, 16'h6586,
// 16'h6663, 16'h6534, 16'h61f6, 16'h5cb8,
// 16'h55a2, 16'h4cc4, 16'h4264, 16'h36a0,
// 16'h29c9, 16'h1c16, 16'h0dd2, 16'hff44,
// 16'hf0bf, 16'he281, 16'hd4e6, 16'hc823,
// 16'hbc83, 16'hb245, 16'ha996, 16'ha2a9,
// 16'h9da2, 16'h9a94, 16'h999c, 16'h9aaf,
// 16'h9dd5, 16'ha2f8, 16'ha9f9, 16'hb2c1,
// 16'hbd0f, 16'hc8c1, 16'hd58c, 16'he339,
// 16'hf173, 16'h2004, 16'h0e86, 16'h1ccc,
// 16'h2a71, 16'h3741, 16'h42ef, 16'h4d41,
// 16'h5606, 16'h5d08, 16'h622b, 16'h6550,
// 16'h6666, 16'h6569, 16'h6261, 16'h5d55,
// 16'h566a, 16'h4dbd, 16'h437a, 16'h37df,
// 16'h2b1a, 16'h1d7e, 16'h0f42, 16'h20bc,
// 16'hf22d, 16'he3ec, 16'hd636, 16'hc95e,
// 16'hbd9f, 16'hb33a, 16'haa60, 16'ha347,
// 16'h9e09, 16'h9acd, 16'h999b, 16'h9a7e,
// 16'h9d6d, 16'ha25e, 16'ha931, 16'hb1cc,
// 16'hbbf7, 16'hc789, 16'hd43a, 16'he1d0,
// 16'hf006, 16'hfe88, 16'h0d1b, 16'h1b60,
// 16'h291f, 16'h3602, 16'h41d6, 16'h4c47,
// 16'h553c, 16'h5c67, 16'h61c0, 16'h6517,
// 16'h6661, 16'h659b, 16'h62c7, 16'h5dea,
// 16'h5734, 16'h4ea8, 16'h4498, 16'h3910,
// 16'h2c72, 16'h1edd, 16'h10b7, 16'h022e,
// 16'hf3a3, 16'he550, 16'hd790, 16'hca98,
// 16'hbec0, 16'hb430, 16'hab31, 16'ha3e7,
// 16'h9e79, 16'h9b09, 16'h99a2, 16'h9a4d,
// 16'h9d0d, 16'ha1c5, 16'ha872, 16'hb0da,
// 16'hbae4, 16'hc651, 16'hd2e9, 16'he06d,
// 16'hee95, 16'hfd13, 16'h0ba9, 16'h19f6,
// 16'h27c9, 16'h34c3, 16'h40b4, 16'h4b50,
// 16'h5466, 16'h5bc8, 16'h614b, 16'h64da,
// 16'h6656, 16'h65ca, 16'h6322, 16'h5e82,
// 16'h57f1, 16'h4f99, 16'h45a7, 16'h3a49,
// 16'h2dbe, 16'h2043, 16'h1226, 16'h03a3,
// 16'hf517, 16'he6b9, 16'hd8e7, 16'hcbdb,
// 16'hbfde, 16'hb530, 16'hac03, 16'ha48c,
// 16'h9eef, 16'h9b48, 16'h99af, 16'h9a25,
// 16'h9cac, 16'ha13b, 16'ha7ad, 16'haff3,
// 16'hb9d0, 16'hc51e, 16'hd19c, 16'hdf0b,
// 16'hed24, 16'hfba0, 16'h0a32, 16'h188f,
// 16'h266e, 16'h3383, 16'h3f90, 16'h4a51,
// 16'h5391, 16'h5b1f, 16'h60d5, 16'h6495,
// 16'h664b, 16'h65ed, 16'h637e, 16'h5f10,
// 16'h58ac, 16'h5086, 16'h46b3, 16'h3b7d,
// 16'h2f09, 16'h21a7, 16'h1393, 16'h0519,
// 16'hf68a, 16'he824, 16'hda42, 16'hcd1c,
// 16'hc104, 16'hb630, 16'hacdc, 16'ha536,
// 16'h9f69, 16'h9b8d, 16'h99c1, 16'h9a20,
// 16'h9c57, 16'ha0ac, 16'ha6f6, 16'haf09,
// 16'hb8c3, 16'hc3ef, 16'hd04f, 16'hddaa,
// 16'hebb7, 16'hfa28, 16'h08c1, 16'h1723,
// 16'h2512, 16'h3242, 16'h3e66, 16'h494f,
// 16'h52b7, 16'h5a73, 16'h6059, 16'h644c,
// 16'h6636, 16'h660f, 16'h63d5, 16'h5f96,
// 16'h5966, 16'h5169, 16'h47c1, 16'h3cac,
// 16'h3051, 16'h230a, 16'h14fd, 16'h0693,
// 16'hf7f9, 16'he994, 16'hdb9b, 16'hce64,
// 16'hc22b, 16'hb735, 16'hadb7, 16'ha5e7,
// 16'h9fe5, 16'h9bdc, 16'h99d5, 16'h99e1,
// 16'h9c05, 16'ha025, 16'ha641, 16'hae26,
// 16'hb7b9, 16'hc2c1, 16'hcf07, 16'hdc4b,
// 16'hea47, 16'hf8b8, 16'h0748, 16'h15b9,
// 16'h23b5, 16'h30f9, 16'h3d3f, 16'h4847,
// 16'h51d9, 16'h59c1, 16'h5fda, 16'h63fc,
// 16'h661e, 16'h662a, 16'h6426, 16'h601a,
// 16'h5a19, 16'h524a, 16'h48c9, 16'h3dd6,
// 16'h319c, 16'h2465, 16'h166c, 16'h0807,
// 16'hf96d, 16'heb02, 16'hdcf8, 16'hcfac,
// 16'hc357, 16'hb83d, 16'hae98, 16'ha69b,
// 16'ha066, 16'h9c2f, 16'h99ef, 16'h99cb,
// 16'h9bb4, 16'h9fa6, 16'ha58d, 16'had4b,
// 16'hb6af, 16'hc19b, 16'hcdbc, 16'hdaf2,
// 16'he8d8, 16'hf744, 16'h05d4, 16'h144b,
// 16'h2255, 16'h2fb2, 16'h3c0f, 16'h4740,
// 16'h50f4, 16'h590c, 16'h5f52, 16'h63ab,
// 16'h65fe, 16'h6642, 16'h646f, 16'h609c,
// 16'h5ac5, 16'h5329, 16'h49cb, 16'h3f20,
// 16'h32e2, 16'h25be, 16'h17de, 16'h0973,
// 16'hfaea, 16'hec6a, 16'hde5b, 16'hd0f6,
// 16'hc485, 16'hb949, 16'haf7f, 16'ha74f,
// 16'ha0f5, 16'h9c7f, 16'h9a13, 16'h99b7,
// 16'h9b69, 16'h9f2d, 16'ha4df, 16'hac6f,
// 16'hb5b1, 16'hc06d, 16'hcc81, 16'hd98d,
// 16'he775, 16'hf5cb, 16'h0461, 16'h12dc,
// 16'h20f5, 16'h2e65, 16'h3ae1, 16'h462f,
// 16'h5010, 16'h5850, 16'h5ec8, 16'h6352,
// 16'h65da, 16'h6654, 16'h64b6, 16'h6111,
// 16'h5b75, 16'h53fb, 16'h4ad3, 16'h401f,
// 16'h3426, 16'h271a, 16'h1945, 16'h0aeb,
// 16'hfc5c, 16'hedda, 16'hdfbe, 16'hd241,
// 16'hc5b7, 16'hba5b, 16'hb064, 16'ha811,
// 16'ha17e, 16'h9cdd, 16'h9a38, 16'h99a9,
// 16'h9b25, 16'h9eb7, 16'ha436, 16'hab9b,
// 16'hb4af, 16'hbf4f, 16'hcb39, 16'hd83b,
// 16'he604, 16'hf45d, 16'h02e9, 16'h116f,
// 16'h1f90, 16'h2d17, 16'h39b0, 16'h451b,
// 16'h4f26, 16'h5791, 16'h5e36, 16'h62f8,
// 16'h65af, 16'h665f, 16'h64f9, 16'h6183,
// 16'h5c1e, 16'h54cb, 16'h4bd3, 16'h413e,
// 16'h3569, 16'h286f, 16'h1ab1, 16'h0c5d,
// 16'hfdd1, 16'hef4b, 16'he120, 16'hd391,
// 16'hc6ec, 16'hbb6d, 16'hb153, 16'ha8d0,
// 16'ha212, 16'h9d3d, 16'h9a62, 16'h99a0,
// 16'h9ae9, 16'h9e41, 16'ha398, 16'haac5,
// 16'hb3b7, 16'hbe2c, 16'hc9fd, 16'hd6e2,
// 16'he49e, 16'hf2e9, 16'h0173, 16'h0ffe,
// 16'h1e2c, 16'h2bc8, 16'h3878, 16'h4408,
// 16'h4e35, 16'h56cc, 16'h5da5, 16'h6291,
// 16'h6584, 16'h6664, 16'h6534, 16'h61f6,
// 16'h5cb9, 16'h55a1, 16'h4cc4, 16'h4264,
// 16'h36a0, 16'h29ca, 16'h1c14, 16'h0dd3,
// 16'hff45, 16'hf0bc, 16'he284, 16'hd4e4,
// 16'hc823, 16'hbc84, 16'hb245, 16'ha994,
// 16'ha2ac, 16'h9d9f, 16'h9a97, 16'h9998,
// 16'h9ab4, 16'h9dd1, 16'ha2fa, 16'ha9f9,
// 16'hb2c0, 16'hbd0f, 16'hc8c3, 16'hd589,
// 16'he33b, 16'hf174, 16'h2020, 16'h0e8a,
// 16'h1cca, 16'h2a72, 16'h3740, 16'h42f0,
// 16'h4d40, 16'h5607, 16'h5d08, 16'h622b,
// 16'h6550, 16'h6666, 16'h656a, 16'h625f,
// 16'h5d57, 16'h5669, 16'h4dbd, 16'h437a,
// 16'h37df, 16'h2b1b, 16'h1d7d, 16'h0f43,
// 16'h20b9, 16'hf231, 16'he3e8, 16'hd63b,
// 16'hc95b, 16'hbda0, 16'hb338, 16'haa62,
// 16'ha344, 16'h9e0e, 16'h9ac9, 16'h999d,
// 16'h9a7c, 16'h9d6e, 16'ha25c, 16'ha935,
// 16'hb1c8, 16'hbbfb, 16'hc785, 16'hd43c,
// 16'he1cf, 16'hf007, 16'hfe89, 16'h0d19,
// 16'h1b61, 16'h291e, 16'h3605, 16'h41d1,
// 16'h4c4d, 16'h5535, 16'h5c6e, 16'h61bb,
// 16'h6519, 16'h6661, 16'h659b, 16'h62c5,
// 16'h5dec, 16'h5732, 16'h4eac, 16'h4493,
// 16'h3915, 16'h2c6c, 16'h1ee4, 16'h10b1,
// 16'h0233, 16'hf39f, 16'he553, 16'hd78e,
// 16'hca99, 16'hbec0, 16'hb430, 16'hab31,
// 16'ha3e7, 16'h9e78, 16'h9b0b, 16'h99a0,
// 16'h9a4e, 16'h9d0e, 16'ha1c3, 16'ha876,
// 16'hb0d5, 16'hbae8, 16'hc64e, 16'hd2eb,
// 16'he06d, 16'hee94, 16'hfd15, 16'h0ba5,
// 16'h19fb, 16'h27c3, 16'h34ca, 16'h40ae,
// 16'h4b53, 16'h5466, 16'h5bc6, 16'h614e,
// 16'h64d7, 16'h6659, 16'h65c8, 16'h6323,
// 16'h5e81, 16'h57f1, 16'h4f9b, 16'h45a5,
// 16'h3a4a, 16'h2dbd, 16'h2044, 16'h1225,
// 16'h03a4, 16'hf516, 16'he6ba, 16'hd8e6,
// 16'hcbdb, 16'hbfde, 16'hb530, 16'hac04,
// 16'ha48b, 16'h9eef, 16'h9b4a, 16'h99ab,
// 16'h9a29, 16'h9caa, 16'ha13b, 16'ha7ae,
// 16'haff3, 16'hb9ce, 16'hc522, 16'hd197,
// 16'hdf0f, 16'hed21, 16'hfba1, 16'h0a32,
// 16'h1890, 16'h266c, 16'h3386, 16'h3f8c,
// 16'h4a54, 16'h538f, 16'h5b20, 16'h60d6,
// 16'h6494, 16'h664a, 16'h65ee, 16'h637e,
// 16'h5f0f, 16'h58ad, 16'h5084, 16'h46b6,
// 16'h3b7a, 16'h2f0c, 16'h21a3, 16'h1396,
// 16'h0519, 16'hf688, 16'he827, 16'hda3f,
// 16'hcd1e, 16'hc104, 16'hb62f, 16'hacdd,
// 16'ha535, 16'h9f69, 16'h9b8f, 16'h99be,
// 16'h9a04, 16'h9c51, 16'ha0b2, 16'ha6f1,
// 16'haf0d, 16'hb8c1, 16'hc3ef, 16'hd04f,
// 16'hddab, 16'hebb5, 16'hfa2b, 16'h08bf,
// 16'h1722, 16'h2515, 16'h323d, 16'h3e6b,
// 16'h494e, 16'h52b5, 16'h5a76, 16'h6055,
// 16'h6450, 16'h6633, 16'h6611, 16'h63d4,
// 16'h5f96, 16'h5967, 16'h5167, 16'h47c4,
// 16'h3ca8, 16'h3055, 16'h2306, 16'h1520,
// 16'h0692, 16'hf7f9, 16'he995, 16'hdb99,
// 16'hce66, 16'hc229, 16'hb737, 16'hadb6,
// 16'ha5e7, 16'h9fe6, 16'h9bda, 16'h99d6,
// 16'h99e3, 16'h9c01, 16'ha029, 16'ha63e,
// 16'hae27, 16'hb7b9, 16'hc2c2, 16'hcf04,
// 16'hdc4e, 16'hea46, 16'hf8b7, 16'h0749,
// 16'h15b9, 16'h23b4, 16'h30fb, 16'h3d3c,
// 16'h484a, 16'h51d6, 16'h59c5, 16'h5fd4,
// 16'h6402, 16'h661a, 16'h662c, 16'h6426,
// 16'h6018, 16'h5a1c, 16'h5248, 16'h48ca,
// 16'h3dd7, 16'h319a, 16'h2466, 16'h166e,
// 16'h0802, 16'hf973, 16'heafd, 16'hdcfc,
// 16'hcfaa, 16'hc357, 16'hb83e, 16'hae97,
// 16'ha69b, 16'ha069, 16'h9c2b, 16'h99f2,
// 16'h99c9, 16'h9bb4, 16'h9fa7, 16'ha58e,
// 16'had47, 16'hb6b4, 16'hc196, 16'hcdc1,
// 16'hdaee, 16'he8db, 16'hf742, 16'h05d5,
// 16'h144b, 16'h2256, 16'h2fb0, 16'h3c12,
// 16'h473d, 16'h50f5, 16'h590d, 16'h5f51,
// 16'h63ab, 16'h65ff, 16'h6640, 16'h6472,
// 16'h6098, 16'h5ac8, 16'h5326, 16'h49cf,
// 16'h3efe, 16'h32e0, 16'h25c3, 16'h17d7,
// 16'h097b, 16'hfae2, 16'hec71, 16'hde56,
// 16'hd0fa, 16'hc482, 16'hb94b, 16'haf7d,
// 16'ha751, 16'ha0f4, 16'h9c7f, 16'h9a14,
// 16'h99b5, 16'h9b6c, 16'h9f2a, 16'ha4e1,
// 16'hac6f, 16'hb5af, 16'hc071, 16'hcc7c,
// 16'hd992, 16'he771, 16'hf5cd, 16'h0462,
// 16'h12d9, 16'h20f8, 16'h2e62, 16'h3ae4,
// 16'h462e, 16'h500f, 16'h5850, 16'h5ec9,
// 16'h6350, 16'h65de, 16'h664f, 16'h64b9,
// 16'h6111, 16'h5b74, 16'h53fb, 16'h4ad3,
// 16'h401f, 16'h3427, 16'h271a, 16'h1943,
// 16'h0aee, 16'hfc59, 16'heddd, 16'hdfbb,
// 16'hd243, 16'hc5b7, 16'hba59, 16'hb067,
// 16'ha80e, 16'ha17f, 16'h9cde, 16'h9a36,
// 16'h99a9, 16'h9b27, 16'h9eb5, 16'ha437,
// 16'hab9b, 16'hb4af, 16'hbf4d, 16'hcb3c,
// 16'hd839, 16'he606, 16'hf45b, 16'h02eb,
// 16'h116b, 16'h1f95, 16'h2d14, 16'h39b0,
// 16'h451d, 16'h4f24, 16'h5792, 16'h5e35,
// 16'h62f9, 16'h65ad, 16'h6662, 16'h64f6,
// 16'h6185, 16'h5c1c, 16'h54ce, 16'h4bce,
// 16'h4144, 16'h3563, 16'h2875, 16'h1aab,
// 16'h0c62, 16'hfdcd, 16'hef4e, 16'he11e,
// 16'hd393, 16'hc6ea, 16'hbb6f, 16'hb151,
// 16'ha8d1, 16'ha213, 16'h9d3a, 16'h9a66,
// 16'h999d, 16'h9aeb, 16'h9e3f, 16'ha399,
// 16'haac4, 16'hb3b9, 16'hbe2a, 16'hc9ff,
// 16'hd6e0, 16'he49f, 16'hf2e7, 16'h0176,
// 16'h0ffb, 16'h1e30, 16'h2bc5, 16'h3878,
// 16'h4409, 16'h4e34, 16'h56cd, 16'h5da5,
// 16'h6290, 16'h6585, 16'h6664, 16'h6533,
// 16'h61f6, 16'h5cba, 16'h559f, 16'h4cc8,
// 16'h425f, 16'h36a5, 16'h29c5, 16'h1c19,
// 16'h0dcf, 16'hff47, 16'hf0bb, 16'he286,
// 16'hd4e1, 16'hc826, 16'hbc83, 16'hb243,
// 16'ha998, 16'ha2a9, 16'h9da0, 16'h9a97,
// 16'h9999, 16'h9ab1, 16'h9dd6, 16'ha2f6,
// 16'ha9fb, 16'hb2be, 16'hbd12, 16'hc8bf,
// 16'hd58f, 16'he335, 16'hf177, 16'h2020,
// 16'h0e89, 16'h1ccb, 16'h2a71, 16'h3742,
// 16'h42ec, 16'h4d45, 16'h5603, 16'h5d0a,
// 16'h622b, 16'h654e, 16'h6668, 16'h6568,
// 16'h6262, 16'h5d54, 16'h566c, 16'h4dba,
// 16'h437c, 16'h37de, 16'h2b1a, 16'h1d80,
// 16'h0f3f, 16'h20be, 16'hf22c, 16'he3ed,
// 16'hd635, 16'hc960, 16'hbd9d, 16'hb33a,
// 16'haa62, 16'ha344, 16'h9e0c, 16'h9acc,
// 16'h999a, 16'h9a7f, 16'h9d6b, 16'ha260,
// 16'ha931, 16'hb1cb, 16'hbbf8, 16'hc788,
// 16'hd43a, 16'he1d2, 16'hf004, 16'hfe8a,
// 16'h0d19, 16'h1b62, 16'h291d, 16'h3605,
// 16'h41d2, 16'h4c4a, 16'h5539, 16'h5c6a,
// 16'h61bf, 16'h6516, 16'h6662, 16'h659b,
// 16'h62c4, 16'h5def, 16'h572e, 16'h4eaf,
// 16'h4492, 16'h3915, 16'h2c6d, 16'h1ee1,
// 16'h10b4, 16'h0231, 16'hf3a1, 16'he552,
// 16'hd78e, 16'hca98, 16'hbec2, 16'hb42e,
// 16'hab33, 16'ha3e5, 16'h9e7a, 16'h9b09,
// 16'h99a1, 16'h9a4f, 16'h9d0a, 16'ha1c9,
// 16'ha86f, 16'hb0dc, 16'hbae2, 16'hc652,
// 16'hd2e9, 16'he06e, 16'hee94, 16'hfd14,
// 16'h0ba6, 16'h19fa, 16'h27c5, 16'h34c8,
// 16'h40b0, 16'h4b51, 16'h5466, 16'h5bc8,
// 16'h614c, 16'h64d8, 16'h665a, 16'h65c4,
// 16'h6329, 16'h5e7c, 16'h57f4, 16'h4f99,
// 16'h45a6, 16'h3a4b, 16'h2dbb, 16'h2047,
// 16'h1220, 16'h03aa, 16'hf510, 16'he6bf,
// 16'hd8e3, 16'hcbdd, 16'hbfdd, 16'hb531,
// 16'hac01, 16'ha48f, 16'h9eec, 16'h9b4b,
// 16'h99ad, 16'h9a25, 16'h9cad, 16'ha13a,
// 16'ha7ad, 16'haff4, 16'hb9cf, 16'hc51f,
// 16'hd19b, 16'hdf0b, 16'hed24, 16'hfba1,
// 16'h0a31, 16'h1890, 16'h266d, 16'h3384,
// 16'h3f90, 16'h4a50, 16'h5392, 16'h5b1e,
// 16'h60d8, 16'h6491, 16'h664e, 16'h65ea,
// 16'h6382, 16'h5f0d, 16'h58ad, 16'h5085,
// 16'h46b4, 16'h3b7d, 16'h2f09, 16'h21a6,
// 16'h1394, 16'h051a, 16'hf688, 16'he826,
// 16'hda3f, 16'hcd1f, 16'hc103, 16'hb630,
// 16'hacdc, 16'ha535, 16'h9f69, 16'h9b90,
// 16'h99bd, 16'h9a03, 16'h9c54, 16'ha0ad,
// 16'ha6f9, 16'haf05, 16'hb8c7, 16'hc3eb,
// 16'hd051, 16'hddab, 16'hebb5, 16'hfa2a,
// 16'h08c0, 16'h1722, 16'h2514, 16'h3240,
// 16'h3e66, 16'h4952, 16'h52b3, 16'h5a77,
// 16'h6055, 16'h644f, 16'h6634, 16'h6610,
// 16'h63d6, 16'h5f93, 16'h596b, 16'h5163,
// 16'h47c7, 16'h3ca5, 16'h3058, 16'h2304,
// 16'h1502, 16'h068f, 16'hf7fd, 16'he990,
// 16'hdb9f, 16'hce60, 16'hc22d, 16'hb736,
// 16'hadb6, 16'ha5e7, 16'h9fe6, 16'h9bda,
// 16'h99d6, 16'h99e3, 16'h9c01, 16'ha029,
// 16'ha63e, 16'hae27, 16'hb7ba, 16'hc2bf,
// 16'hcf08, 16'hdc4b, 16'hea47, 16'hf8b8,
// 16'h0748, 16'h15b9, 16'h23b5, 16'h30f9,
// 16'h3d3f, 16'h4848, 16'h51d7, 16'h59c3,
// 16'h5fd7, 16'h63ff, 16'h661d, 16'h662a,
// 16'h6425, 16'h601a, 16'h5a1a, 16'h524a,
// 16'h48ca, 16'h3dd5, 16'h319b, 16'h2467,
// 16'h166b, 16'h0807, 16'hf96e, 16'heb20,
// 16'hdcfa, 16'hcfab, 16'hc357, 16'hb83d,
// 16'hae98, 16'ha69a, 16'ha069, 16'h9c2b,
// 16'h99f3, 16'h99c7, 16'h9bb8, 16'h9fa3,
// 16'ha590, 16'had46, 16'hb6b6, 16'hc193,
// 16'hcdc5, 16'hdae9, 16'he8df, 16'hf740,
// 16'h05d5, 16'h144c, 16'h2254, 16'h2fb2,
// 16'h3c11, 16'h473d, 16'h50f6, 16'h590c,
// 16'h5f51, 16'h63ad, 16'h65fd, 16'h6642,
// 16'h6470, 16'h6099, 16'h5ac8, 16'h5326,
// 16'h49cf, 16'h3efd, 16'h32e3, 16'h25be,
// 16'h17db, 16'h0979, 16'hfae3, 16'hec71,
// 16'hde56, 16'hd0f8, 16'hc485, 16'hb949,
// 16'haf7e, 16'ha751, 16'ha0f3, 16'h9c80,
// 16'h9a14, 16'h99b3, 16'h9b6f, 16'h9f28,
// 16'ha4e1, 16'hac71, 16'hb5ac, 16'hc073,
// 16'hcc7b, 16'hd992, 16'he773, 16'hf5cb,
// 16'h0463, 16'h12d9, 16'h20f7, 16'h2e64,
// 16'h3ae1, 16'h4631, 16'h500e, 16'h5850,
// 16'h5ec8, 16'h6352, 16'h65da, 16'h6655,
// 16'h64b3, 16'h6115, 16'h5b72, 16'h53fd,
// 16'h4ad1, 16'h4020, 16'h3427, 16'h2719,
// 16'h1945, 16'h0aec, 16'hfc5a, 16'heddd,
// 16'hdfbb, 16'hd242, 16'hc5b8, 16'hba59,
// 16'hb067, 16'ha80e, 16'ha180, 16'h9cda,
// 16'h9a3b, 16'h99a6, 16'h9b29, 16'h9eb3,
// 16'ha438, 16'hab9a, 16'hb4b0, 16'hbf4e,
// 16'hcb3a, 16'hd839, 16'he607, 16'hf45b,
// 16'h02eb, 16'h116b, 16'h1f94, 16'h2d14,
// 16'h39b3, 16'h4518, 16'h4f29, 16'h578d,
// 16'h5e3a, 16'h62f5, 16'h65b1, 16'h665f,
// 16'h64f7, 16'h6186, 16'h5c1a, 16'h54d0,
// 16'h4bce, 16'h4142, 16'h3566, 16'h2871,
// 16'h1aaf, 16'h0c5f, 16'hfdcf, 16'hef4d,
// 16'he11d, 16'hd394, 16'hc6ea, 16'hbb70,
// 16'hb14f, 16'ha8d3, 16'ha210, 16'h9d3e,
// 16'h9a63, 16'h99a0, 16'h9ae6, 16'h9e46,
// 16'ha392, 16'haacb, 16'hb3b2, 16'hbe30,
// 16'hc9fb, 16'hd6e2, 16'he4a0, 16'hf2e4,
// 16'h0179, 16'h0ffa, 16'h1e2e, 16'h2bc8,
// 16'h3876, 16'h440a, 16'h4e34, 16'h56cc,
// 16'h5da6, 16'h628e, 16'h6589, 16'h665f,
// 16'h6538, 16'h61f2, 16'h5cbc, 16'h559f,
// 16'h4cc7, 16'h4261, 16'h36a2, 16'h29c9,
// 16'h1c15, 16'h0dd2, 16'hff45, 16'hf0bc,
// 16'he286, 16'hd4e2, 16'hc823, 16'hbc86,
// 16'hb241, 16'ha99a, 16'ha2a7, 16'h9da1,
// 16'h9a97, 16'h9999, 16'h9ab1, 16'h9dd6,
// 16'ha2f4, 16'ha9fe, 16'hb2bc, 16'hbd14,
// 16'hc8bd, 16'hd58f, 16'he336, 16'hf176,
// 16'h2001, 16'h0e89, 16'h1cc9, 16'h2a73,
// 16'h3741, 16'h42ed, 16'h4d44, 16'h5603,
// 16'h5d0a, 16'h622b, 16'h654e, 16'h6668,
// 16'h6569, 16'h625f, 16'h5d58, 16'h5667,
// 16'h4dbf, 16'h437a, 16'h37dd, 16'h2b1d,
// 16'h1d7b, 16'h0f45, 16'h20b9, 16'hf22f,
// 16'he3eb, 16'hd636, 16'hc960, 16'hbd9c,
// 16'hb33c, 16'haa5e, 16'ha349, 16'h9e08,
// 16'h9ace, 16'h999b, 16'h9a7b, 16'h9d71,
// 16'ha25a, 16'ha935, 16'hb1ca, 16'hbbf8,
// 16'hc787, 16'hd43b, 16'he1d1, 16'hf004,
// 16'hfe8c, 16'h0d16, 16'h1b63, 16'h291f,
// 16'h3601, 16'h41d6, 16'h4c48, 16'h5539,
// 16'h5c6c, 16'h61bb, 16'h651a, 16'h665f,
// 16'h659d, 16'h62c4, 16'h5ded, 16'h5731,
// 16'h4eac, 16'h4494, 16'h3914, 16'h2c6e,
// 16'h1ee1, 16'h10b4, 16'h0230, 16'hf3a2,
// 16'he552, 16'hd78c, 16'hca9e, 16'hbeb9,
// 16'hb436, 16'hab2d, 16'ha3e9, 16'h9e79,
// 16'h9b08, 16'h99a2, 16'h9a4e, 16'h9d0b,
// 16'ha1c9, 16'ha86f, 16'hb0db, 16'hbae3,
// 16'hc652, 16'hd2e9, 16'he06e, 16'hee93,
// 16'hfd15, 16'h0ba7, 16'h19f8, 16'h27c8,
// 16'h34c3, 16'h40b5, 16'h4b4e, 16'h5468,
// 16'h5bc7, 16'h614c, 16'h64d9, 16'h6657,
// 16'h65ca, 16'h6320, 16'h5e85, 16'h57ed,
// 16'h4f9e, 16'h45a4, 16'h3a4a, 16'h2dbd,
// 16'h2043, 16'h1227, 16'h03a2, 16'hf517,
// 16'he6ba, 16'hd8e6, 16'hcbdb, 16'hbfdf,
// 16'hb52e, 16'hac05, 16'ha48c, 16'h9eed,
// 16'h9b4b, 16'h99ad, 16'h9a25, 16'h9cae,
// 16'ha138, 16'ha7af, 16'haff3, 16'hb9cf,
// 16'hc51f, 16'hd19c, 16'hdf09, 16'hed27,
// 16'hfb9d, 16'h0a35, 16'h188d, 16'h266f,
// 16'h3383, 16'h3f90, 16'h4a51, 16'h5390,
// 16'h5b20, 16'h60d6, 16'h6493, 16'h664c,
// 16'h65ec, 16'h6380, 16'h5f0e, 16'h58ad,
// 16'h5085, 16'h46b4, 16'h3b7d, 16'h2f08,
// 16'h21a8, 16'h1392, 16'h051b, 16'hf688,
// 16'he825, 16'hda41, 16'hcd1d, 16'hc104,
// 16'hb630, 16'hacdb, 16'ha537, 16'h9f68,
// 16'h9b8f, 16'h99bf, 16'h9a02, 16'h9c54,
// 16'ha0af, 16'ha6f3, 16'haf0d, 16'hb8c0,
// 16'hc3f1, 16'hd04d, 16'hddac, 16'hebb4,
// 16'hfa2d, 16'h08bd, 16'h1724, 16'h2513,
// 16'h323f, 16'h3e6a, 16'h494d, 16'h52b7,
// 16'h5a73, 16'h6059, 16'h644d, 16'h6635,
// 16'h6610, 16'h63d4, 16'h5f96, 16'h5967,
// 16'h5168, 16'h47c2, 16'h3cab, 16'h3052,
// 16'h2308, 16'h1520, 16'h0690, 16'hf7fc,
// 16'he992, 16'hdb9b, 16'hce65, 16'hc22a,
// 16'hb737, 16'hadb6, 16'ha5e6, 16'h9fe6,
// 16'h9bdc, 16'h99d4, 16'h99e5, 16'h9c20,
// 16'ha028, 16'ha640, 16'hae25, 16'hb7bc,
// 16'hc2bf, 16'hcf06, 16'hdc4e, 16'hea44,
// 16'hf8ba, 16'h0747, 16'h15b9, 16'h23b6,
// 16'h30f7, 16'h3d41, 16'h4846, 16'h51d9,
// 16'h59c3, 16'h5fd5, 16'h6401, 16'h661b,
// 16'h662c, 16'h6425, 16'h601a, 16'h5a19,
// 16'h524b, 16'h48c8, 16'h3dd7, 16'h319b,
// 16'h2465, 16'h166e, 16'h0804, 16'hf970,
// 16'heaff, 16'hdcfa, 16'hcfac, 16'hc357,
// 16'hb83c, 16'hae9a, 16'ha697, 16'ha06c,
// 16'h9c2a, 16'h99f2, 16'h99c9, 16'h9bb4,
// 16'h9fa7, 16'ha58d, 16'had4a, 16'hb6b1,
// 16'hc198, 16'hcdbf, 16'hdaf0, 16'he8d9,
// 16'hf745, 16'h05d2, 16'h144d, 16'h2255,
// 16'h2fb0, 16'h3c12, 16'h473d, 16'h50f6,
// 16'h590c, 16'h5f51, 16'h63ab, 16'h65ff,
// 16'h6640, 16'h6472, 16'h6097, 16'h5acb,
// 16'h5323, 16'h49d1, 16'h3efb, 16'h32e4,
// 16'h25be, 16'h17dd, 16'h0976, 16'hfae6,
// 16'hec6d, 16'hde5a, 16'hd0f5, 16'hc488,
// 16'hb946, 16'haf80, 16'ha750, 16'ha0f4,
// 16'h9c7f, 16'h9a14, 16'h99b4, 16'h9b6d,
// 16'h9f2b, 16'ha4df, 16'hac71, 16'hb5ac,
// 16'hc074, 16'hcc7b, 16'hd992, 16'he771,
// 16'hf5ce, 16'h045f, 16'h12de, 16'h20f3,
// 16'h2e66, 16'h3ae1, 16'h462f, 16'h500f,
// 16'h5851, 16'h5ec7, 16'h6352, 16'h65dc,
// 16'h6651, 16'h64b9, 16'h610f, 16'h5b75,
// 16'h53fd, 16'h4ad0, 16'h4022, 16'h3425,
// 16'h2719, 16'h1947, 16'h0ae9, 16'hfc5e,
// 16'hedd8, 16'hdfbf, 16'hd241, 16'hc5b6,
// 16'hba5e, 16'hb060, 16'ha813, 16'ha17e,
// 16'h9cdc, 16'h9a3a, 16'h99a5, 16'h9b2a,
// 16'h9eb2, 16'ha43a, 16'hab99, 16'hb4af,
// 16'hbf4f, 16'hcb3a, 16'hd839, 16'he608,
// 16'hf458, 16'h02ee, 16'h116a, 16'h1f94,
// 16'h2d16, 16'h39ae, 16'h451f, 16'h4f22,
// 16'h5793, 16'h5e36, 16'h62f6, 16'h65b2,
// 16'h665e, 16'h64f7, 16'h6187, 16'h5c19,
// 16'h54cf, 16'h4bd0, 16'h4140, 16'h3568,
// 16'h2870, 16'h1ab0, 16'h0c5d, 16'hfdd1,
// 16'hef4b, 16'he11f, 16'hd393, 16'hc6eb,
// 16'hbb6d, 16'hb153, 16'ha8d0, 16'ha213,
// 16'h9d3b, 16'h9a65, 16'h999e, 16'h9ae9,
// 16'h9e44, 16'ha392, 16'haacb, 16'hb3b4,
// 16'hbe2d, 16'hc9fe, 16'hd6df, 16'he4a1,
// 16'hf2e6, 16'h0176, 16'h0ffc, 16'h1e2e,
// 16'h2bc7, 16'h3877, 16'h4409, 16'h4e34,
// 16'h56cf, 16'h5da1, 16'h6294, 16'h6582,
// 16'h6666, 16'h6533, 16'h61f4, 16'h5cbd,
// 16'h559d, 16'h4cc8, 16'h4261, 16'h36a1,
// 16'h29ca, 16'h1c16, 16'h0dd0, 16'hff46,
// 16'hf0be, 16'he280, 16'hd4e9, 16'hc81e,
// 16'hbc89, 16'hb240, 16'ha999, 16'ha2a7,
// 16'h9da3, 16'h9a95, 16'h999a, 16'h9ab0,
// 16'h9dd6, 16'ha2f5, 16'ha9fe, 16'hb2bb,
// 16'hbd14, 16'hc8bd, 16'hd590, 16'he334,
// 16'hf178, 16'hffff, 16'h0e8a, 16'h1cca,
// 16'h2a72, 16'h3740, 16'h42ef, 16'h4d42,
// 16'h5604, 16'h5d0a, 16'h622b, 16'h654e,
// 16'h6669, 16'h6567, 16'h6261, 16'h5d55,
// 16'h566b, 16'h4dbc, 16'h437c, 16'h37dc,
// 16'h2b1c, 16'h1d7d, 16'h0f43, 16'h20bb,
// 16'hf22e, 16'he3eb, 16'hd636, 16'hc960,
// 16'hbd9c, 16'hb33d, 16'haa5d, 16'ha348,
// 16'h9e0a, 16'h9acc, 16'h999c, 16'h9a7d,
// 16'h9d6c, 16'ha25f, 16'ha931, 16'hb1cc,
// 16'hbbf9, 16'hc785, 16'hd43d, 16'he1cf,
// 16'hf005, 16'hfe8b, 16'h0d18, 16'h1b62,
// 16'h291e, 16'h3603, 16'h41d3, 16'h4c4b,
// 16'h5538, 16'h5c6b, 16'h61be, 16'h6516,
// 16'h6663, 16'h6599, 16'h62c8, 16'h5deb,
// 16'h5732, 16'h4eab, 16'h4493, 16'h3916,
// 16'h2c6d, 16'h1ee2, 16'h10b2, 16'h0232,
// 16'hf3a0, 16'he553, 16'hd78e, 16'hca99,
// 16'hbec0, 16'hb430, 16'hab31, 16'ha3e6,
// 16'h9e7a, 16'h9b09, 16'h99a1, 16'h9a4f,
// 16'h9d0a, 16'ha1c9, 16'ha86f, 16'hb0dc,
// 16'hbae2, 16'hc651, 16'hd2eb, 16'he06d,
// 16'hee93, 16'hfd17, 16'h0ba2, 16'h19fd,
// 16'h27c4, 16'h34c7, 16'h40b2, 16'h4b50,
// 16'h5467, 16'h5bc6, 16'h614e, 16'h64d6,
// 16'h665b, 16'h65c6, 16'h6324, 16'h5e82,
// 16'h57ee, 16'h4f9d, 16'h45a4, 16'h3a4b,
// 16'h2dbc, 16'h2046, 16'h1221, 16'h03a9,
// 16'hf511, 16'he6bd, 16'hd8e6, 16'hcbda,
// 16'hbfe0, 16'hb52f, 16'hac02, 16'ha48e,
// 16'h9eee, 16'h9b48, 16'h99b0, 16'h9a23,
// 16'h9caf, 16'ha137, 16'ha7b1, 16'haff0,
// 16'hb9d2, 16'hc51d, 16'hd19c, 16'hdf0b,
// 16'hed25, 16'hfb9e, 16'h0a35, 16'h188c,
// 16'h2672, 16'h337f, 16'h3f94, 16'h4a4c,
// 16'h5396, 16'h5b1b, 16'h60d9, 16'h6491,
// 16'h664d, 16'h65ec, 16'h6380, 16'h5f0d,
// 16'h58af, 16'h5082, 16'h46b8, 16'h3b79,
// 16'h2f0b, 16'h21a6, 16'h1393, 16'h051b,
// 16'hf687, 16'he827, 16'hda3f, 16'hcd1e,
// 16'hc104, 16'hb630, 16'hacdb, 16'ha536,
// 16'h9f69, 16'h9b8f, 16'h99bf, 16'h9a01,
// 16'h9c56, 16'ha0ab, 16'ha6f9, 16'haf07,
// 16'hb8c4, 16'hc3ef, 16'hd04d, 16'hddae,
// 16'hebb2, 16'hfa2e, 16'h08bb, 16'h1727,
// 16'h2511, 16'h3240, 16'h3e69, 16'h494d,
// 16'h52b8, 16'h5a73, 16'h6057, 16'h644f,
// 16'h6634, 16'h6610, 16'h63d4, 16'h5f96,
// 16'h5968, 16'h5166, 16'h47c5, 16'h3ca6,
// 16'h3057, 16'h2305, 16'h1502, 16'h068f,
// 16'hf7fc, 16'he992, 16'hdb9b, 16'hce66,
// 16'hc228, 16'hb738, 16'hadb5, 16'ha5e8,
// 16'h9fe4, 16'h9bdd, 16'h99d2, 16'h99e7,
// 16'h9bfe, 16'ha02b, 16'ha63d, 16'hae27,
// 16'hb7ba, 16'hc2bf, 16'hcf0a, 16'hdc47,
// 16'hea4c, 16'hf8b3, 16'h074b, 16'h15b9,
// 16'h23b3, 16'h30fb, 16'h3d3f, 16'h4845,
// 16'h51dc, 16'h59bf, 16'h5fda, 16'h63fd,
// 16'h661d, 16'h662b, 16'h6426, 16'h6018,
// 16'h5a1d, 16'h5245, 16'h48ce, 16'h3dd2,
// 16'h31a0, 16'h2460, 16'h1672, 16'h0820,
// 16'hf974, 16'heafc, 16'hdcfc, 16'hcfaa,
// 16'hc359, 16'hb83a, 16'hae9b, 16'ha698,
// 16'ha06a, 16'h9c2c, 16'h99f0, 16'h99cb,
// 16'h9bb3, 16'h9fa8, 16'ha58c, 16'had4b,
// 16'hb6b0, 16'hc199, 16'hcdbf, 16'hdaef,
// 16'he8db, 16'hf742, 16'h05d5, 16'h144b,
// 16'h2256, 16'h2fb0, 16'h3c12, 16'h473d,
// 16'h50f6, 16'h590b, 16'h5f53, 16'h63ab,
// 16'h65fe, 16'h6642, 16'h646f, 16'h609a,
// 16'h5ac8, 16'h5325, 16'h49d1, 16'h3efa,
// 16'h32e5, 16'h25bd, 16'h17dc, 16'h0977,
// 16'hfae7, 16'hec6a, 16'hde5d, 16'hd0f4,
// 16'hc486, 16'hb949, 16'haf7e, 16'ha750,
// 16'ha0f4, 16'h9c80, 16'h9a13, 16'h99b5,
// 16'h9b6d, 16'h9f28, 16'ha4e3, 16'hac6d,
// 16'hb5b1, 16'hc06f, 16'hcc7d, 16'hd993,
// 16'he76f, 16'hf5d0, 16'h045e, 16'h12dd,
// 16'h20f5, 16'h2e64, 16'h3ae3, 16'h462d,
// 16'h5012, 16'h584d, 16'h5ecb, 16'h634f,
// 16'h65de, 16'h6650, 16'h64b8, 16'h6112,
// 16'h5b73, 16'h53fc, 16'h4ad3, 16'h401f,
// 16'h3426, 16'h271b, 16'h1943, 16'h0aed,
// 16'hfc5b, 16'hedda, 16'hdfbe, 16'hd241,
// 16'hc5b8, 16'hba58, 16'hb068, 16'ha80d,
// 16'ha181, 16'h9cdb, 16'h9a39, 16'h99a7,
// 16'h9b29, 16'h9eb2, 16'ha43a, 16'hab99,
// 16'hb4af, 16'hbf4f, 16'hcb39, 16'hd83c,
// 16'he603, 16'hf45e, 16'h02e8, 16'h116e,
// 16'h1f93, 16'h2d14, 16'h39b2, 16'h451b,
// 16'h4f25, 16'h5791, 16'h5e36, 16'h62f8,
// 16'h65af, 16'h6661, 16'h64f5, 16'h6187,
// 16'h5c1b, 16'h54cd, 16'h4bd1, 16'h4141,
// 16'h3566, 16'h2871, 16'h1ab1, 16'h0c5b,
// 16'hfdd3, 16'hef4a, 16'he120, 16'hd392,
// 16'hc6eb, 16'hbb6e, 16'hb151, 16'ha8d3,
// 16'ha210, 16'h9d3c, 16'h9a66, 16'h999c,
// 16'h9aeb, 16'h9e42, 16'ha394, 16'haaca,
// 16'hb3b3, 16'hbe30, 16'hc9f9, 16'hd6e6,
// 16'he49a, 16'hf2eb, 16'h0173, 16'h0ffd,
// 16'h1e2f, 16'h2bc4, 16'h387c, 16'h4404,
// 16'h4e37, 16'h56cd, 16'h5da3, 16'h6293,
// 16'h6583, 16'h6664, 16'h6534, 16'h61f6,
// 16'h5cb9, 16'h55a1, 16'h4cc5, 16'h4262,
// 16'h36a2, 16'h29c8, 16'h1c18, 16'h0dcf,
// 16'hff46, 16'hf0bd, 16'he282, 16'hd4e8,
// 16'hc81f, 16'hbc87, 16'hb242, 16'ha998,
// 16'ha2a8, 16'h9da2, 16'h9a95, 16'h999b,
// 16'h9ab0, 16'h9dd5, 16'ha2f7, 16'ha9fa,
// 16'hb2c1, 16'hbd0e, 16'hc8c3, 16'hd58b,
// 16'he337, 16'hf178, 16'hfffd, 16'h0e8e,
// 16'h1cc6, 16'h2a74, 16'h3740, 16'h42ee,
// 16'h4d43, 16'h5604, 16'h5d0a, 16'h622a,
// 16'h6550, 16'h6667, 16'h6568, 16'h6261,
// 16'h5d56, 16'h5669, 16'h4dbf, 16'h4378,
// 16'h37e0, 16'h2b19, 16'h1d80, 16'h0f40,
// 16'h20bc, 16'hf230, 16'he3e6, 16'hd63d,
// 16'hc959, 16'hbda2, 16'hb338, 16'haa60,
// 16'ha347, 16'h9e0a, 16'h9acd, 16'h999b,
// 16'h9a7c, 16'h9d6e, 16'ha25d, 16'ha933,
// 16'hb1ca, 16'hbbf9, 16'hc787, 16'hd439,
// 16'he1d4, 16'hf001, 16'hfe8e, 16'h0d16,
// 16'h1b62, 16'h291f, 16'h3603, 16'h41d2,
// 16'h4c4e, 16'h5533, 16'h5c70, 16'h61b9,
// 16'h651a, 16'h6660, 16'h659d, 16'h62c3,
// 16'h5def, 16'h572e, 16'h4eaf, 16'h4492,
// 16'h3914, 16'h2c6f, 16'h1ee0, 16'h10b5,
// 16'h022f, 16'hf3a3, 16'he550, 16'hd78f,
// 16'hca9b, 16'hbebc, 16'hb433, 16'hab31,
// 16'ha3e4, 16'h9e7e, 16'h9b04, 16'h99a5,
// 16'h9a4c, 16'h9d0d, 16'ha1c7, 16'ha870,
// 16'hb0da, 16'hbae5, 16'hc64f, 16'hd2ec,
// 16'he06b, 16'hee96, 16'hfd12, 16'h0ba9,
// 16'h19f7, 16'h27c8, 16'h34c5, 16'h40b1,
// 16'h4b53, 16'h5463, 16'h5bcb, 16'h6149,
// 16'h64db, 16'h6657, 16'h65c7, 16'h6325,
// 16'h5e80, 16'h57f2, 16'h4f99, 16'h45a7,
// 16'h3a49, 16'h2dbe, 16'h2043, 16'h1225,
// 16'h03a5, 16'hf514, 16'he6bc, 16'hd8e5,
// 16'hcbdb, 16'hbfe0, 16'hb52c, 16'hac07,
// 16'ha48a, 16'h9ef0, 16'h9b48, 16'h99ad,
// 16'h9a27, 16'h9cad, 16'ha138, 16'ha7b1,
// 16'hafee, 16'hb9d4, 16'hc51d, 16'hd19b,
// 16'hdf0c, 16'hed23, 16'hfba1, 16'h0a31,
// 16'h1890, 16'h266e, 16'h3382, 16'h3f93,
// 16'h4a4c, 16'h5396, 16'h5b1b, 16'h60d8,
// 16'h6493, 16'h664d, 16'h65ea, 16'h6382,
// 16'h5f0b, 16'h58b1, 16'h5081, 16'h46b8,
// 16'h3b79, 16'h2f0b, 16'h21a6, 16'h1393,
// 16'h051b, 16'hf687, 16'he827, 16'hda3e,
// 16'hcd21, 16'hc101, 16'hb631, 16'hacdb,
// 16'ha537, 16'h9f67, 16'h9b91, 16'h99bd,
// 16'h9a03, 16'h9c54, 16'ha0ae, 16'ha6f5,
// 16'haf0a, 16'hb8c4, 16'hc3eb, 16'hd054,
// 16'hdda6, 16'hebb9, 16'hfa29, 16'h08bf,
// 16'h1724, 16'h2512, 16'h3240, 16'h3e68,
// 16'h4950, 16'h52b4, 16'h5a76, 16'h6056,
// 16'h644f, 16'h6634, 16'h6610, 16'h63d4,
// 16'h5f97, 16'h5966, 16'h5169, 16'h47c2,
// 16'h3ca9, 16'h3055, 16'h2306, 16'h1520,
// 16'h0692, 16'hf7f9, 16'he994, 16'hdb9b,
// 16'hce63, 16'hc22c, 16'hb735, 16'hadb8,
// 16'ha5e5, 16'h9fe7, 16'h9bd9, 16'h99d8,
// 16'h99e0, 16'h9c05, 16'ha025, 16'ha640,
// 16'hae27, 16'hb7b9, 16'hc2c0, 16'hcf08,
// 16'hdc4a, 16'hea48, 16'hf8b7, 16'h0749,
// 16'h15b9, 16'h23b4, 16'h30fa, 16'h3d3f,
// 16'h4846, 16'h51da, 16'h59c1, 16'h5fd8,
// 16'h63ff, 16'h661b, 16'h662c, 16'h6425,
// 16'h601a, 16'h5a1a, 16'h5248, 16'h48cc,
// 16'h3dd4, 16'h319c, 16'h2466, 16'h166b,
// 16'h0808, 16'hf96d, 16'heb01, 16'hdcfa,
// 16'hcfa9, 16'hc35a, 16'hb83a, 16'hae9c,
// 16'ha696, 16'ha06d, 16'h9c27, 16'h99f5,
// 16'h99c7, 16'h9bb7, 16'h9fa4, 16'ha590,
// 16'had45, 16'hb6b6, 16'hc195, 16'hcdc1,
// 16'hdaed, 16'he8dd, 16'hf740, 16'h05d7,
// 16'h1449, 16'h2256, 16'h2fb0, 16'h3c13,
// 16'h473c, 16'h50f7, 16'h5909, 16'h5f55,
// 16'h63a8, 16'h6602, 16'h663e, 16'h6473,
// 16'h6097, 16'h5ac9, 16'h5326, 16'h49cf,
// 16'h3efd, 16'h32e3, 16'h25be, 16'h17dc,
// 16'h0977, 16'hfae6, 16'hec6c, 16'hde5c,
// 16'hd0f2, 16'hc48a, 16'hb945, 16'haf80,
// 16'ha751, 16'ha0f1, 16'h9c83, 16'h9a11,
// 16'h99b6, 16'h9b6c, 16'h9f2a, 16'ha4e1,
// 16'hac70, 16'hb5ad, 16'hc072, 16'hcc7b,
// 16'hd994, 16'he770, 16'hf5ce, 16'h045f,
// 16'h12dc, 16'h20f7, 16'h2e62, 16'h3ae4,
// 16'h462d, 16'h5010, 16'h5850, 16'h5ec9,
// 16'h6350, 16'h65dd, 16'h6651, 16'h64b7,
// 16'h6113, 16'h5b71, 16'h53ff, 16'h4ad0,
// 16'h4021, 16'h3425, 16'h271b, 16'h1943,
// 16'h0aed, 16'hfc5b, 16'hedda, 16'hdfbd,
// 16'hd243, 16'hc5b5, 16'hba5d, 16'hb062,
// 16'ha812, 16'ha17c, 16'h9ce1, 16'h9a33,
// 16'h99ac, 16'h9b25, 16'h9eb4, 16'ha43a,
// 16'hab98, 16'hb4b1, 16'hbf4c, 16'hcb3c,
// 16'hd838, 16'he608, 16'hf459, 16'h02ed,
// 16'h1169, 16'h1f96, 16'h2d14, 16'h39b0,
// 16'h451c, 16'h4f26, 16'h578f, 16'h5e3a,
// 16'h62f3, 16'h65b3, 16'h665d, 16'h64fa,
// 16'h6182, 16'h5c1e, 16'h54cd, 16'h4bcf,
// 16'h4143, 16'h3564, 16'h2873, 16'h1aaf,
// 16'h0c5c, 16'hfdd3, 16'hef49, 16'he122,
// 16'hd38f, 16'hc6ee, 16'hbb6c, 16'hb152,
// 16'ha8d3, 16'ha20e, 16'h9d41, 16'h9a5f,
// 16'h99a3, 16'h9ae6, 16'h9e45, 16'ha392,
// 16'haaca, 16'hb3b5, 16'hbe2d, 16'hc9fd,
// 16'hd6e1, 16'he49e, 16'hf2e9, 16'h0174,
// 16'h0ffc, 16'h1e30, 16'h2bc3, 16'h387c,
// 16'h4405, 16'h4e37, 16'h56cc, 16'h5da4,
// 16'h6291, 16'h6585, 16'h6664, 16'h6533,
// 16'h61f6, 16'h5cbb, 16'h559d, 16'h4cca,
// 16'h425d, 16'h36a6, 16'h29c7, 16'h1c16,
// 16'h0dd1, 16'hff45, 16'hf0be, 16'he283,
// 16'hd4e4, 16'hc823, 16'hbc84, 16'hb245,
// 16'ha994, 16'ha2ad, 16'h9d9d, 16'h9a99,
// 16'h9997, 16'h9ab4, 16'h9dd2, 16'ha2f9,
// 16'ha9f9, 16'hb2c0, 16'hbd11, 16'hc8c0,
// 16'hd58c, 16'he338, 16'hf176, 16'hffff,
// 16'h0e8c, 16'h1cc6, 16'h2a77, 16'h373b,
// 16'h42f4, 16'h4d3d, 16'h5609, 16'h5d06,
// 16'h622d, 16'h654e, 16'h6668, 16'h6567,
// 16'h6263, 16'h5d53, 16'h566d, 16'h4dba,
// 16'h437c, 16'h37dd, 16'h2b1c, 16'h1d7c,
// 16'h0f45, 16'h20b8, 16'hf230, 16'he3ea,
// 16'hd637, 16'hc95e, 16'hbd9f, 16'hb339,
// 16'haa61, 16'ha346, 16'h9e09, 16'h9ace,
// 16'h999b, 16'h9a7d, 16'h9d6d, 16'ha25e,
// 16'ha932, 16'hb1cb, 16'hbbf9, 16'hc786,
// 16'hd43c, 16'he1d0, 16'hf005, 16'hfe8a,
// 16'h0d19, 16'h1b62, 16'h291c, 16'h3606,
// 16'h41d1, 16'h4c4d, 16'h5536, 16'h5c6c,
// 16'h61bd, 16'h6516, 16'h6664, 16'h659a,
// 16'h62c5, 16'h5dee, 16'h572f, 16'h4ead,
// 16'h4494, 16'h3913, 16'h2c6f, 16'h1ee2,
// 16'h10b2, 16'h0232, 16'hf39f, 16'he554,
// 16'hd78d, 16'hca9b, 16'hbebd, 16'hb432,
// 16'hab31, 16'ha3e4, 16'h9e7e, 16'h9b03,
// 16'h99a8, 16'h9a49, 16'h9d0e, 16'ha1c7,
// 16'ha86f, 16'hb0dd, 16'hbae2, 16'hc651,
// 16'hd2eb, 16'he06b, 16'hee96, 16'hfd14,
// 16'h0ba6, 16'h19f9, 16'h27c7, 16'h34c4,
// 16'h40b5, 16'h4b4e, 16'h5468, 16'h5bc6,
// 16'h614c, 16'h64da, 16'h6657, 16'h65c8,
// 16'h6324, 16'h5e80, 16'h57f2, 16'h4f99,
// 16'h45a7, 16'h3a48, 16'h2dbf, 16'h2043,
// 16'h1225, 16'h03a5, 16'hf514, 16'he6bc,
// 16'hd8e6, 16'hcbd9, 16'hbfe2, 16'hb52b,
// 16'hac08, 16'ha488, 16'h9ef1, 16'h9b48,
// 16'h99ae, 16'h9a24, 16'h9caf, 16'ha137,
// 16'ha7b1, 16'haff1, 16'hb9d0, 16'hc51f,
// 16'hd19b, 16'hdf0b, 16'hed25, 16'hfb9f,
// 16'h0a32, 16'h1890, 16'h266e, 16'h3383,
// 16'h3f90, 16'h4a4f, 16'h5393, 16'h5b1f,
// 16'h60d4, 16'h6497, 16'h6647, 16'h65f1,
// 16'h637c, 16'h5f10, 16'h58ad, 16'h5083,
// 16'h46b8, 16'h3b78, 16'h2f0e, 16'h21a2,
// 16'h1396, 16'h0519, 16'hf688, 16'he827,
// 16'hda40, 16'hcd1c, 16'hc105, 16'hb630,
// 16'hacda, 16'ha539, 16'h9f65, 16'h9b91,
// 16'h99bf, 16'h9a20, 16'h9c57, 16'ha0ac,
// 16'ha6f6, 16'haf09, 16'hb8c3, 16'hc3ef,
// 16'hd050, 16'hdda9, 16'hebb7, 16'hfa29,
// 16'h08c0, 16'h1724, 16'h2511, 16'h3242,
// 16'h3e67, 16'h494f, 16'h52b7, 16'h5a72,
// 16'h6059, 16'h644e, 16'h6633, 16'h6612,
// 16'h63d2, 16'h5f99, 16'h5964, 16'h516a,
// 16'h47c1, 16'h3ca9, 16'h3057, 16'h2302,
// 16'h1506, 16'h068b, 16'hf7ff, 16'he991,
// 16'hdb9a, 16'hce66, 16'hc22a, 16'hb736,
// 16'hadb7, 16'ha5e6, 16'h9fe5, 16'h9bdd,
// 16'h99d3, 16'h99e6, 16'h9bfe, 16'ha02c,
// 16'ha63b, 16'hae2a, 16'hb7b8, 16'hc2c0,
// 16'hcf08, 16'hdc4b, 16'hea47, 16'hf8b8,
// 16'h0747, 16'h15bb, 16'h23b3, 16'h30fa,
// 16'h3d40, 16'h4845, 16'h51db, 16'h59c0,
// 16'h5fd9, 16'h63fd, 16'h661f, 16'h6628,
// 16'h6428, 16'h6017, 16'h5a1d, 16'h5247,
// 16'h48cb, 16'h3dd5, 16'h319c, 16'h2464,
// 16'h1670, 16'h0801, 16'hf974, 16'heafb,
// 16'hdcfd, 16'hcfa9, 16'hc359, 16'hb83d,
// 16'hae97, 16'ha69b, 16'ha067, 16'h9c2e,
// 16'h99f0, 16'h99ca, 16'h9bb5, 16'h9fa5,
// 16'ha58f, 16'had47, 16'hb6b4, 16'hc195,
// 16'hcdc3, 16'hdaeb, 16'he8dd, 16'hf743,
// 16'h05d1, 16'h1450, 16'h2250, 16'h2fb6,
// 16'h3c0d, 16'h4741, 16'h50f2, 16'h590f,
// 16'h5f4f, 16'h63ad, 16'h65fe, 16'h6640,
// 16'h6473, 16'h6095, 16'h5acc, 16'h5322,
// 16'h49d3, 16'h3ef9, 16'h32e6, 16'h25bc,
// 16'h17dd, 16'h0977, 16'hfae6, 16'hec6c,
// 16'hde5b, 16'hd0f5, 16'hc487, 16'hb948,
// 16'haf7e, 16'ha751, 16'ha0f3, 16'h9c81,
// 16'h9a12, 16'h99b6, 16'h9b6c, 16'h9f2a,
// 16'ha4e1, 16'hac6e, 16'hb5b0, 16'hc071,
// 16'hcc7c, 16'hd992, 16'he771, 16'hf5cd,
// 16'h0461, 16'h12dc, 16'h20f4, 16'h2e66,
// 16'h3ae0, 16'h4631, 16'h500d, 16'h5853,
// 16'h5ec4, 16'h6356, 16'h65d8, 16'h6654,
// 16'h64b6, 16'h6113, 16'h5b71, 16'h5420,
// 16'h4ace, 16'h4023, 16'h3425, 16'h2719,
// 16'h1945, 16'h0aee, 16'hfc57, 16'hede0,
// 16'hdfb7, 16'hd247, 16'hc5b4, 16'hba5c,
// 16'hb064, 16'ha80f, 16'ha181, 16'h9cda,
// 16'h9a3b, 16'h99a5, 16'h9b2a, 16'h9eb1,
// 16'ha43c, 16'hab96, 16'hb4b3, 16'hbf4b,
// 16'hcb3c, 16'hd839, 16'he607, 16'hf45b,
// 16'h02e9, 16'h116e, 16'h1f91, 16'h2d18,
// 16'h39af, 16'h451c, 16'h4f25, 16'h5790,
// 16'h5e38, 16'h62f6, 16'h65b1, 16'h665e,
// 16'h64f8, 16'h6186, 16'h5c1a, 16'h54cf,
// 16'h4bcf, 16'h4141, 16'h3567, 16'h2872,
// 16'h1aad, 16'h0c61, 16'hfdcd, 16'hef4f,
// 16'he11d, 16'hd393, 16'hc6eb, 16'hbb6e,
// 16'hb152, 16'ha8d1, 16'ha212, 16'h9d3b,
// 16'h9a66, 16'h999d, 16'h9aea, 16'h9e42,
// 16'ha394, 16'haaca, 16'hb3b3, 16'hbe30,
// 16'hc9fa, 16'hd6e3, 16'he49d, 16'hf2ea,
// 16'h0172, 16'h0fff, 16'h1e2c, 16'h2bc7,
// 16'h3879, 16'h4407, 16'h4e35, 16'h56ce,
// 16'h5da3, 16'h6291, 16'h6585, 16'h6663,
// 16'h6536, 16'h61f3, 16'h5cbd, 16'h559b,
// 16'h4ccb, 16'h425e, 16'h36a5, 16'h29c7,
// 16'h1c16, 16'h0dd1, 16'hff45, 16'hf0bf,
// 16'he280, 16'hd4e8, 16'hc820, 16'hbc86,
// 16'hb243, 16'ha996, 16'ha2aa, 16'h9da2,
// 16'h9a94, 16'h999b, 16'h9ab0, 16'h9dd5,
// 16'ha2f7, 16'ha9fb, 16'hb2be, 16'hbd12,
// 16'hc8bf, 16'hd58d, 16'he338, 16'hf175,
// 16'h2001, 16'h0e89, 16'h1cca, 16'h2a72,
// 16'h3741, 16'h42ee, 16'h4d42, 16'h5605,
// 16'h5d09, 16'h622b, 16'h654f, 16'h6667,
// 16'h6569, 16'h6260, 16'h5d57, 16'h5668,
// 16'h4dbe, 16'h437a, 16'h37df, 16'h2b1a,
// 16'h1d7e, 16'h0f41, 16'h20bd, 16'hf22d,
// 16'he3eb, 16'hd637, 16'hc95e, 16'hbd9f,
// 16'hb339, 16'haa61, 16'ha345, 16'h9e0d,
// 16'h9ac9, 16'h999f, 16'h9a7a, 16'h9d6f,
// 16'ha25d, 16'ha933, 16'hb1ca, 16'hbbfa,
// 16'hc784, 16'hd43f, 16'he1cd, 16'hf008,
// 16'hfe87, 16'h0d1b, 16'h1b61, 16'h291d,
// 16'h3606, 16'h41cf, 16'h4c4f, 16'h5534,
// 16'h5c6e, 16'h61bb, 16'h6519, 16'h6661,
// 16'h659a, 16'h62c7, 16'h5deb, 16'h5732,
// 16'h4eac, 16'h4493, 16'h3915, 16'h2c6c,
// 16'h1ee4, 16'h10b1, 16'h0233, 16'hf39e,
// 16'he554, 16'hd78e, 16'hca99, 16'hbec0,
// 16'hb42f, 16'hab31, 16'ha3e8, 16'h9e77,
// 16'h9b0c, 16'h999e, 16'h9a51, 16'h9d0a,
// 16'ha1c8, 16'ha870, 16'hb0db, 16'hbae3,
// 16'hc652, 16'hd2e9, 16'he06d, 16'hee95,
// 16'hfd14, 16'h0ba7, 16'h19f7, 16'h27c8,
// 16'h34c6, 16'h40b1, 16'h4b52, 16'h5463,
// 16'h5bcb, 16'h614a, 16'h64da, 16'h6657,
// 16'h65c8, 16'h6324, 16'h5e80, 16'h57f2,
// 16'h4f99, 16'h45a8, 16'h3a48, 16'h2dbe,
// 16'h2043, 16'h1225, 16'h03a5, 16'hf515,
// 16'he6ba, 16'hd8e7, 16'hcbda, 16'hbfdf,
// 16'hb52f, 16'hac03, 16'ha48c, 16'h9ef0,
// 16'h9b47, 16'h99b0, 16'h9a23, 16'h9cae,
// 16'ha13a, 16'ha7ad, 16'haff3, 16'hb9d1,
// 16'hc51c, 16'hd19e, 16'hdf09, 16'hed24,
// 16'hfba3, 16'h0a2e, 16'h1892, 16'h266d,
// 16'h3382, 16'h3f93, 16'h4a4d, 16'h5394,
// 16'h5b1d, 16'h60d6, 16'h6496, 16'h6647,
// 16'h65f2, 16'h637b, 16'h5f10, 16'h58ae,
// 16'h5081, 16'h46ba, 16'h3b77, 16'h2f0e,
// 16'h21a2, 16'h1396, 16'h0518, 16'hf68c,
// 16'he821, 16'hda44, 16'hcd1b, 16'hc105,
// 16'hb630, 16'hacdb, 16'ha537, 16'h9f68,
// 16'h9b8f, 16'h99bf, 16'h9a01, 16'h9c56,
// 16'ha0ad, 16'ha6f5, 16'haf0a, 16'hb8c3,
// 16'hc3ee, 16'hd050, 16'hdda9, 16'hebb7,
// 16'hfa2a, 16'h08bf, 16'h1724, 16'h2512,
// 16'h323f, 16'h3e6b, 16'h494b, 16'h52bb,
// 16'h5a6f, 16'h605b, 16'h644c, 16'h6634,
// 16'h6612, 16'h63d2, 16'h5f98, 16'h5966,
// 16'h5167, 16'h47c4, 16'h3ca7, 16'h3057,
// 16'h2304, 16'h1503, 16'h068e, 16'hf7fd,
// 16'he991, 16'hdb9c, 16'hce65, 16'hc229,
// 16'hb738, 16'hadb4, 16'ha5e9, 16'h9fe4,
// 16'h9bdc, 16'h99d5, 16'h99e2, 16'h9c04,
// 16'ha025, 16'ha642, 16'hae25, 16'hb7ba,
// 16'hc2c0, 16'hcf07, 16'hdc4c, 16'hea47,
// 16'hf8b7, 16'h0749, 16'h15b9, 16'h23b4,
// 16'h30fa, 16'h3d3e, 16'h4848, 16'h51d9,
// 16'h59c0, 16'h5fd9, 16'h63fe, 16'h661c,
// 16'h662d, 16'h6423, 16'h601c, 16'h5a18,
// 16'h524b, 16'h48c9, 16'h3dd5, 16'h319f,
// 16'h2460, 16'h1672, 16'h0801, 16'hf972,
// 16'heaff, 16'hdcfa, 16'hcfaa, 16'hc358,
// 16'hb83e, 16'hae97, 16'ha69b, 16'ha068,
// 16'h9c2d, 16'h99f0, 16'h99ca, 16'h9bb5,
// 16'h9fa5, 16'ha590, 16'had46, 16'hb6b4,
// 16'hc197, 16'hcdbf, 16'hdaf0, 16'he8d9,
// 16'hf744, 16'h05d4, 16'h144a, 16'h2257,
// 16'h2fb0, 16'h3c11, 16'h473e, 16'h50f5,
// 16'h590d, 16'h5f50, 16'h63ae, 16'h65fa,
// 16'h6645, 16'h646f, 16'h6099, 16'h5aca,
// 16'h5322, 16'h49d3, 16'h3efa, 16'h32e4,
// 16'h25c0, 16'h17d9, 16'h0979, 16'hfae5,
// 16'hec6d, 16'hde5b, 16'hd0f5, 16'hc485,
// 16'hb94a, 16'haf7c, 16'ha754, 16'ha0ef,
// 16'h9c85, 16'h9a0f, 16'h99b8, 16'h9b69,
// 16'h9f2d, 16'ha4de, 16'hac73, 16'hb5ac,
// 16'hc071, 16'hcc7d, 16'hd991, 16'he773,
// 16'hf5cc, 16'h0461, 16'h12db, 16'h20f7,
// 16'h2e62, 16'h3ae5, 16'h462b, 16'h5013,
// 16'h584e, 16'h5ec8, 16'h6353, 16'h65da,
// 16'h6653, 16'h64b6, 16'h6112, 16'h5b73,
// 16'h53ff, 16'h4ace, 16'h4023, 16'h3424,
// 16'h271b, 16'h1945, 16'h0aec, 16'hfc5a,
// 16'heddb, 16'hdfbe, 16'hd240, 16'hc5ba,
// 16'hba58, 16'hb065, 16'ha810, 16'ha17e,
// 16'h9cde, 16'h9a37, 16'h99a9, 16'h9b26,
// 16'h9eb5, 16'ha438, 16'hab99, 16'hb4b1,
// 16'hbf4d, 16'hcb3b, 16'hd838, 16'he609,
// 16'hf457, 16'h02ef, 16'h1169, 16'h1f94,
// 16'h2d16, 16'h39af, 16'h451d, 16'h4f25,
// 16'h5790, 16'h5e38, 16'h62f5, 16'h65b2,
// 16'h665e, 16'h64f8, 16'h6186, 16'h5c19,
// 16'h54d1, 16'h4bcd, 16'h4143, 16'h3566,
// 16'h2871, 16'h1aaf, 16'h0c5f, 16'hfdcf,
// 16'hef4e, 16'he11c, 16'hd394, 16'hc6eb,
// 16'hbb6d, 16'hb154, 16'ha8cf, 16'ha212,
// 16'h9d3c, 16'h9a65, 16'h999d, 16'h9aec,
// 16'h9e3f, 16'ha398, 16'haac5, 16'hb3b8,
// 16'hbe2c, 16'hc9fd, 16'hd6e2, 16'he49d,
// 16'hf2e9, 16'h0175, 16'h0ffc, 16'h1e2e,
// 16'h2bc7, 16'h3877, 16'h4409, 16'h4e35,
// 16'h56cc, 16'h5da5, 16'h6291, 16'h6583,
// 16'h6665, 16'h6534, 16'h61f4, 16'h5cbd,
// 16'h559c, 16'h4cc9, 16'h4261, 16'h36a1,
// 16'h29ca, 16'h1c15, 16'h0dd2, 16'hff45,
// 16'hf0bd, 16'he283, 16'hd4e5, 16'hc822,
// 16'hbc85, 16'hb244, 16'ha995, 16'ha2ac,
// 16'h9d9e, 16'h9a98, 16'h9999, 16'h9ab1,
// 16'h9dd4, 16'ha2f9, 16'ha9f8, 16'hb2c2,
// 16'hbd0d, 16'hc8c4, 16'hd58b, 16'he337,
// 16'hf176, 16'h2020, 16'h0e8a, 16'h1ccb,
// 16'h2a70, 16'h3742, 16'h42ed, 16'h4d44,
// 16'h5603, 16'h5d0b, 16'h6229, 16'h6551,
// 16'h6665, 16'h656b, 16'h625f, 16'h5d56,
// 16'h566b, 16'h4dba, 16'h437f, 16'h37da,
// 16'h2b1e, 16'h1d7c, 16'h0f42, 16'h20bc,
// 16'hf22f, 16'he3e9, 16'hd639, 16'hc95c,
// 16'hbda0, 16'hb339, 16'haa61, 16'ha346,
// 16'h9e09, 16'h9acf, 16'h9998, 16'h9a81,
// 16'h9d69, 16'ha262, 16'ha92f, 16'hb1cc,
// 16'hbbf9, 16'hc785, 16'hd43e, 16'he1ce,
// 16'hf007, 16'hfe89, 16'h0d18, 16'h1b63,
// 16'h291d, 16'h3605, 16'h41d2, 16'h4c4b,
// 16'h5538, 16'h5c6b, 16'h61bd, 16'h6518,
// 16'h6661, 16'h659b, 16'h62c6, 16'h5deb,
// 16'h5733, 16'h4eaa, 16'h4495, 16'h3914,
// 16'h2c6e, 16'h1ee1, 16'h10b3, 16'h0232,
// 16'hf3a0, 16'he553, 16'hd78c, 16'hca9c,
// 16'hbebd, 16'hb433, 16'hab2f, 16'ha3e6,
// 16'h9e7b, 16'h9b08, 16'h99a3, 16'h9a4c,
// 16'h9d0d, 16'ha1c6, 16'ha872, 16'hb0da,
// 16'hbae3, 16'hc652, 16'hd2e8, 16'he06f,
// 16'hee92, 16'hfd17, 16'h0ba4, 16'h19fb,
// 16'h27c5, 16'h34c5, 16'h40b4, 16'h4b4e,
// 16'h5469, 16'h5bc5, 16'h614e, 16'h64d7,
// 16'h665a, 16'h65c6, 16'h6325, 16'h5e7f,
// 16'h57f3, 16'h4f99, 16'h45a8, 16'h3a47,
// 16'h2dbf, 16'h2043, 16'h1225, 16'h03a5,
// 16'hf514, 16'he6bc, 16'hd8e5, 16'hcbdc,
// 16'hbfde, 16'hb52e, 16'hac06, 16'ha48a,
// 16'h9ef0, 16'h9b48, 16'h99ae, 16'h9a25,
// 16'h9cae, 16'ha139, 16'ha7af, 16'haff1,
// 16'hb9d1, 16'hc51d, 16'hd19e, 16'hdf08,
// 16'hed27, 16'hfb9d, 16'h0a35, 16'h188d,
// 16'h266f, 16'h3383, 16'h3f90, 16'h4a51,
// 16'h5390, 16'h5b20, 16'h60d6, 16'h6494,
// 16'h664a, 16'h65ee, 16'h637e, 16'h5f10,
// 16'h58ab, 16'h5086, 16'h46b3, 16'h3b7e,
// 16'h2f08, 16'h21a7, 16'h1392, 16'h051b,
// 16'hf688, 16'he825, 16'hda41, 16'hcd1d,
// 16'hc105, 16'hb62e, 16'hacdd, 16'ha535,
// 16'h9f6a, 16'h9b8e, 16'h99bf, 16'h9a02,
// 16'h9c54, 16'ha0af, 16'ha6f4, 16'haf0a,
// 16'hb8c4, 16'hc3ed, 16'hd050, 16'hddaa,
// 16'hebb6, 16'hfa2b, 16'h08bf, 16'h1722,
// 16'h2514, 16'h323f, 16'h3e6a, 16'h494d,
// 16'h52b7, 16'h5a73, 16'h6059, 16'h644d,
// 16'h6634, 16'h6611, 16'h63d3, 16'h5f98,
// 16'h5965, 16'h5169, 16'h47c1, 16'h3cab,
// 16'h3052, 16'h2309, 16'h14ff, 16'h0691,
// 16'hf7fb, 16'he992, 16'hdb9c, 16'hce64,
// 16'hc22b, 16'hb735, 16'hadb9, 16'ha5e3,
// 16'h9fe9, 16'h9bd9, 16'h99d6, 16'h99e3,
// 16'h9c02, 16'ha027, 16'ha641, 16'hae24,
// 16'hb7bc, 16'hc2bf, 16'hcf08, 16'hdc4a,
// 16'hea49, 16'hf8b5, 16'h074c, 16'h15b6,
// 16'h23b6, 16'h30f9, 16'h3d3f, 16'h4848,
// 16'h51d8, 16'h59c1, 16'h5fd9, 16'h63fe,
// 16'h661d, 16'h662b, 16'h6425, 16'h6019,
// 16'h5a1c, 16'h5247, 16'h48cc, 16'h3dd4,
// 16'h319c, 16'h2466, 16'h166b, 16'h0808,
// 16'hf96c, 16'heb04, 16'hdcf5, 16'hcfaf,
// 16'hc355, 16'hb83e, 16'hae99, 16'ha698,
// 16'ha06b, 16'h9c2b, 16'h99f0, 16'h99cb,
// 16'h9bb4, 16'h9fa6, 16'ha58e, 16'had49,
// 16'hb6b2, 16'hc197, 16'hcdc0, 16'hdaed,
// 16'he8de, 16'hf73f, 16'h05d8, 16'h1447,
// 16'h2259, 16'h2fad, 16'h3c15, 16'h473a,
// 16'h50f9, 16'h5909, 16'h5f53, 16'h63ab,
// 16'h65fe, 16'h6642, 16'h6470, 16'h6099,
// 16'h5ac8, 16'h5326, 16'h49cf, 16'h3efc,
// 16'h32e4, 16'h25be, 16'h17db, 16'h0978,
// 16'hfae5, 16'hec6e, 16'hde5a, 16'hd0f4,
// 16'hc488, 16'hb947, 16'haf7f, 16'ha751,
// 16'ha0f2, 16'h9c82, 16'h9a12, 16'h99b4,
// 16'h9b6f, 16'h9f26, 16'ha4e5, 16'hac6d,
// 16'hb5af, 16'hc071, 16'hcc7d, 16'hd990,
// 16'he774, 16'hf5ca, 16'h0465, 16'h12d7,
// 16'h20f9, 16'h2e61, 16'h3ae4, 16'h462f,
// 16'h500e, 16'h5852, 16'h5ec6, 16'h6353,
// 16'h65dc, 16'h6650, 16'h64b9, 16'h6110,
// 16'h5b75, 16'h53fb, 16'h4ad4, 16'h401c,
// 16'h342b, 16'h2716, 16'h1946, 16'h0aec,
// 16'hfc59, 16'heddf, 16'hdfb9, 16'hd244,
// 16'hc5b6, 16'hba5a, 16'hb066, 16'ha80f,
// 16'ha17f, 16'h9cdc, 16'h9a39, 16'h99a7,
// 16'h9b28, 16'h9eb4, 16'ha439, 16'hab97,
// 16'hb4b4, 16'hbf49, 16'hcb3f, 16'hd836,
// 16'he609, 16'hf459, 16'h02ec, 16'h116b,
// 16'h1f94, 16'h2d15, 16'h39b1, 16'h451a,
// 16'h4f27, 16'h578f, 16'h5e39, 16'h62f5,
// 16'h65b1, 16'h665f, 16'h64f7, 16'h6186,
// 16'h5c1a, 16'h54cf, 16'h4bd0, 16'h4140,
// 16'h3567, 16'h2872, 16'h1aac, 16'h0c63,
// 16'hfdcb, 16'hef4f, 16'he11e, 16'hd392,
// 16'hc6ec, 16'hbb6d, 16'hb152, 16'ha8d2,
// 16'ha211, 16'h9d3b, 16'h9a67, 16'h999b,
// 16'h9aec, 16'h9e41, 16'ha395, 16'haac9,
// 16'hb3b4, 16'hbe2e, 16'hc9fc, 16'hd6e3,
// 16'he49c, 16'hf2ea, 16'h0174, 16'h0ffc,
// 16'h1e30, 16'h2bc3, 16'h387c, 16'h4405,
// 16'h4e37, 16'h56cc, 16'h5da3, 16'h6294,
// 16'h6581, 16'h6666, 16'h6533, 16'h61f5,
// 16'h5cbb, 16'h559f, 16'h4cc6, 16'h4263,
// 16'h36a0, 16'h29cb, 16'h1c14, 16'h0dd2,
// 16'hff46, 16'hf0bc, 16'he285, 16'hd4e2,
// 16'hc825, 16'hbc83, 16'hb245, 16'ha996,
// 16'ha2a9, 16'h9da1, 16'h9a97, 16'h9997,
// 16'h9ab5, 16'h9dd0, 16'ha2fb, 16'ha9f8,
// 16'hb2c1, 16'hbd0e, 16'hc8c4, 16'hd588,
// 16'he33c, 16'hf173, 16'h2020, 16'h0e8c,
// 16'h1cc6, 16'h2a77, 16'h373d, 16'h42ef,
// 16'h4d43, 16'h5603, 16'h5d0c, 16'h6228,
// 16'h6551, 16'h6666, 16'h656a, 16'h625f,
// 16'h5d57, 16'h5669, 16'h4dbd, 16'h437b,
// 16'h37dd, 16'h2b1c, 16'h1d7d, 16'h0f42,
// 16'h20bc, 16'hf22e, 16'he3e9, 16'hd63a,
// 16'hc95b, 16'hbda2, 16'hb336, 16'haa63,
// 16'ha344, 16'h9e0c, 16'h9acc, 16'h999b,
// 16'h9a7e, 16'h9d6b, 16'ha25f, 16'ha932,
// 16'hb1cb, 16'hbbfa, 16'hc784, 16'hd43d,
// 16'he1cf, 16'hf007, 16'hfe88, 16'h0d1a,
// 16'h1b61, 16'h291e, 16'h3605, 16'h41d1,
// 16'h4c4b, 16'h5539, 16'h5c69, 16'h61c1,
// 16'h6513, 16'h6665, 16'h6598, 16'h62c7,
// 16'h5dec, 16'h5731, 16'h4ead, 16'h4492,
// 16'h3915, 16'h2c6e, 16'h1ee1, 16'h10b4,
// 16'h0230, 16'hf3a2, 16'he551, 16'hd790,
// 16'hca98, 16'hbebf, 16'hb431, 16'hab32,
// 16'ha3e4, 16'h9e7c, 16'h9b08, 16'h99a0,
// 16'h9a51, 16'h9d08, 16'ha1ca, 16'ha86f,
// 16'hb0db, 16'hbae4, 16'hc64f, 16'hd2ec,
// 16'he06b, 16'hee97, 16'hfd12, 16'h0ba8,
// 16'h19f7, 16'h27c8, 16'h34c6, 16'h40b1,
// 16'h4b52, 16'h5464, 16'h5bca, 16'h614a,
// 16'h64da, 16'h6657, 16'h65c9, 16'h6323,
// 16'h5e81, 16'h57f0, 16'h4f9b, 16'h45a6,
// 16'h3a4a, 16'h2dbc, 16'h2045, 16'h1224,
// 16'h03a5, 16'hf515, 16'he6ba, 16'hd8e7,
// 16'hcbdb, 16'hbfde, 16'hb52f, 16'hac04,
// 16'ha48d, 16'h9eee, 16'h9b48, 16'h99af,
// 16'h9a24, 16'h9caf, 16'ha138, 16'ha7af,
// 16'haff2, 16'hb9d0, 16'hc51e, 16'hd19d,
// 16'hdf09, 16'hed25, 16'hfba0, 16'h0a32,
// 16'h188f, 16'h266e, 16'h3383, 16'h3f91,
// 16'h4a4f, 16'h5393, 16'h5b1d, 16'h60d8,
// 16'h6492, 16'h664d, 16'h65eb, 16'h6381,
// 16'h5f0d, 16'h58ae, 16'h5083, 16'h46b8,
// 16'h3b78, 16'h2f0d, 16'h21a3, 16'h1396,
// 16'h0518, 16'hf68b, 16'he822, 16'hda44,
// 16'hcd1a, 16'hc106, 16'hb62f, 16'hacdc,
// 16'ha536, 16'h9f68, 16'h9b8f, 16'h99bf,
// 16'h9a02, 16'h9c55, 16'ha0ad, 16'ha6f6,
// 16'haf08, 16'hb8c6, 16'hc3eb, 16'hd053,
// 16'hdda7, 16'hebb8, 16'hfa29, 16'h08c0,
// 16'h1723, 16'h2514, 16'h323d, 16'h3e6c,
// 16'h494b, 16'h52ba, 16'h5a71, 16'h6059,
// 16'h644d, 16'h6636, 16'h660e, 16'h63d6,
// 16'h5f95, 16'h5967, 16'h5168, 16'h47c3,
// 16'h3ca8, 16'h3055, 16'h2307, 16'h14ff,
// 16'h0692, 16'hf7fa, 16'he993, 16'hdb9b,
// 16'hce65, 16'hc229, 16'hb738, 16'hadb5,
// 16'ha5e7, 16'h9fe6, 16'h9bdb, 16'h99d4,
// 16'h99e5, 16'h9c20, 16'ha028, 16'ha641,
// 16'hae23, 16'hb7bd, 16'hc2bd, 16'hcf0a,
// 16'hdc49, 16'hea49, 16'hf8b5, 16'h074b,
// 16'h15b7, 16'h23b6, 16'h30f8, 16'h3d41,
// 16'h4844, 16'h51dd, 16'h59bd, 16'h5fdb,
// 16'h63fe, 16'h661b, 16'h662d, 16'h6423,
// 16'h601c, 16'h5a19, 16'h5249, 16'h48cb,
// 16'h3dd3, 16'h319f, 16'h2462, 16'h1670,
// 16'h0802, 16'hf972, 16'heafd, 16'hdcfc,
// 16'hcfab, 16'hc355, 16'hb840, 16'hae96,
// 16'ha69a, 16'ha06b, 16'h9c29, 16'h99f4,
// 16'h99c7, 16'h9bb6, 16'h9fa6, 16'ha58d,
// 16'had4a, 16'hb6b1, 16'hc199, 16'hcdbd,
// 16'hdaf1, 16'he8d9, 16'hf744, 16'h05d5,
// 16'h1448, 16'h225a, 16'h2fab, 16'h3c18,
// 16'h4737, 16'h50fa, 16'h590a, 16'h5f52,
// 16'h63ac, 16'h65fd, 16'h6641, 16'h6472,
// 16'h6097, 16'h5acb, 16'h5323, 16'h49d1,
// 16'h3efb, 16'h32e3, 16'h25c1, 16'h17d9,
// 16'h0979, 16'hfae5, 16'hec6b, 16'hde5e,
// 16'hd0f1, 16'hc48b, 16'hb944, 16'haf81,
// 16'ha74f, 16'ha0f4, 16'h9c80, 16'h9a14,
// 16'h99b4, 16'h9b6c, 16'h9f2b, 16'ha4df,
// 16'hac72, 16'hb5ad, 16'hc071, 16'hcc7c,
// 16'hd992, 16'he772, 16'hf5cd, 16'h0461,
// 16'h12da, 16'h20f7, 16'h2e63, 16'h3ae3,
// 16'h462f, 16'h500f, 16'h5850, 16'h5ec7,
// 16'h6354, 16'h65d9, 16'h6655, 16'h64b3,
// 16'h6115, 16'h5b72, 16'h53fe, 16'h4acf,
// 16'h4022, 16'h3425, 16'h271b, 16'h1944,
// 16'h0aeb, 16'hfc5c, 16'hedda, 16'hdfbd,
// 16'hd243, 16'hc5b5, 16'hba5c, 16'hb064,
// 16'ha80f, 16'ha182, 16'h9cd7, 16'h9a3e,
// 16'h99a3, 16'h9b2b, 16'h9eb2, 16'ha439,
// 16'hab99, 16'hb4b1, 16'hbf4c, 16'hcb3d,
// 16'hd837, 16'he608, 16'hf45a, 16'h02eb,
// 16'h116c, 16'h1f94, 16'h2d14, 16'h39b1,
// 16'h451c, 16'h4f25, 16'h5791, 16'h5e37,
// 16'h62f5, 16'h65b3, 16'h665c, 16'h64fa,
// 16'h6185, 16'h5c18, 16'h54d4, 16'h4bc8,
// 16'h4149, 16'h3560, 16'h2876, 16'h1aab,
// 16'h0c62, 16'hfdcd, 16'hef4f, 16'he11c,
// 16'hd394, 16'hc6ea, 16'hbb6f, 16'hb151,
// 16'ha8d2, 16'ha211, 16'h9d3c, 16'h9a65,
// 16'h999d, 16'h9aeb, 16'h9e41, 16'ha396,
// 16'haac7, 16'hb3b7, 16'hbe2c, 16'hc9fd,
// 16'hd6e1, 16'he49f, 16'hf2e7, 16'h0177,
// 16'h0ff9, 16'h1e31, 16'h2bc4, 16'h387a,
// 16'h4407, 16'h4e35, 16'h56cd, 16'h5da4,
// 16'h6291, 16'h6585, 16'h6663, 16'h6534,
// 16'h61f6, 16'h5cba, 16'h55a0, 16'h4cc5,
// 16'h4263, 16'h36a1, 16'h29ca, 16'h1c14,
// 16'h0dd3, 16'hff43, 16'hf0c0, 16'he282,
// 16'hd4e3, 16'hc824, 16'hbc83, 16'hb245,
// 16'ha997, 16'ha2a8, 16'h9da2, 16'h9a94,
// 16'h999c, 16'h9aaf, 16'h9dd7, 16'ha2f6,
// 16'ha9fa, 16'hb2bf, 16'hbd11, 16'hc8c1,
// 16'hd58c, 16'he338, 16'hf174, 16'h2002,
// 16'h0e88, 16'h1ccb, 16'h2a71, 16'h3742,
// 16'h42ed, 16'h4d42, 16'h5606, 16'h5d08,
// 16'h622c, 16'h654f, 16'h6665, 16'h656d,
// 16'h625b, 16'h5d5c, 16'h5664, 16'h4dc1,
// 16'h4378, 16'h37e0, 16'h2b1a, 16'h1d7e,
// 16'h0f41, 16'h20bd, 16'hf22d, 16'he3ec,
// 16'hd636, 16'hc95e, 16'hbd9f, 16'hb339,
// 16'haa62, 16'ha344, 16'h9e0c, 16'h9acb,
// 16'h999c, 16'h9a7d, 16'h9d6d, 16'ha25e,
// 16'ha932, 16'hb1cb, 16'hbbf8, 16'hc787,
// 16'hd43c, 16'he1cf, 16'hf007, 16'hfe87,
// 16'h0d1c, 16'h1b5e, 16'h2922, 16'h3620,
// 16'h41d6, 16'h4c48, 16'h5539, 16'h5c6b,
// 16'h61bd, 16'h6518, 16'h6661, 16'h659b,
// 16'h62c6, 16'h5deb, 16'h5733, 16'h4eaa,
// 16'h4495, 16'h3914, 16'h2c6d, 16'h1ee3,
// 16'h10b1, 16'h0234, 16'hf39d, 16'he556,
// 16'hd78a, 16'hca9d, 16'hbebd, 16'hb431,
// 16'hab32, 16'ha3e4, 16'h9e7c, 16'h9b07,
// 16'h99a2, 16'h9a4f, 16'h9d0a, 16'ha1c9,
// 16'ha86f, 16'hb0db, 16'hbae4, 16'hc650,
// 16'hd2eb, 16'he06c, 16'hee95, 16'hfd15,
// 16'h0ba4, 16'h19fb, 16'h27c6, 16'h34c5,
// 16'h40b4, 16'h4b4d, 16'h546a, 16'h5bc4,
// 16'h6150, 16'h64d5, 16'h665b, 16'h65c5,
// 16'h6326, 16'h5e7f, 16'h57f2, 16'h4f9a,
// 16'h45a6, 16'h3a49, 16'h2dbe, 16'h2043,
// 16'h1225, 16'h03a5, 16'hf514, 16'he6bd,
// 16'hd8e4, 16'hcbdc, 16'hbfdd, 16'hb531,
// 16'hac02, 16'ha48f, 16'h9eeb, 16'h9b4c,
// 16'h99aa, 16'h9a29, 16'h9cac, 16'ha139,
// 16'ha7af, 16'haff1, 16'hb9d2, 16'hc51d,
// 16'hd19c, 16'hdf0b, 16'hed23, 16'hfba2,
// 16'h0a31, 16'h188f, 16'h266f, 16'h3381,
// 16'h3f93, 16'h4a4d, 16'h5395, 16'h5b1c,
// 16'h60d7, 16'h6495, 16'h6648, 16'h65f0,
// 16'h637d, 16'h5f0f, 16'h58ad, 16'h5084,
// 16'h46b6, 16'h3b7a, 16'h2f0c, 16'h21a3,
// 16'h1396, 16'h0519, 16'hf689, 16'he825,
// 16'hda40, 16'hcd1e, 16'hc104, 16'hb630,
// 16'hacdc, 16'ha535, 16'h9f68, 16'h9b90,
// 16'h99bf, 16'h9a02, 16'h9c54, 16'ha0ae,
// 16'ha6f4, 16'haf0c, 16'hb8c2, 16'hc3ed,
// 16'hd052, 16'hdda8, 16'hebb7, 16'hfa2b,
// 16'h08bc, 16'h1728, 16'h250e, 16'h3244,
// 16'h3e65, 16'h4951, 16'h52b5, 16'h5a73,
// 16'h605a, 16'h644c, 16'h6635, 16'h6610,
// 16'h63d3, 16'h5f99, 16'h5964, 16'h516a,
// 16'h47c1, 16'h3ca9, 16'h3056, 16'h2305,
// 16'h1502, 16'h068e, 16'hf7fe, 16'he98f,
// 16'hdb9f, 16'hce62, 16'hc22b, 16'hb736,
// 16'hadb7, 16'ha5e5, 16'h9fe8, 16'h9bd8,
// 16'h99d9, 16'h99e0, 16'h9c04, 16'ha026,
// 16'ha63f, 16'hae28, 16'hb7b9, 16'hc2c0,
// 16'hcf08, 16'hdc49, 16'hea4a, 16'hf8b5,
// 16'h074a, 16'h15b9, 16'h23b3, 16'h30fc,
// 16'h3d3c, 16'h484a, 16'h51d7, 16'h59c3,
// 16'h5fd7, 16'h63fe, 16'h661e, 16'h6629,
// 16'h6428, 16'h6017, 16'h5a1c, 16'h5247,
// 16'h48cd, 16'h3dd2, 16'h319f, 16'h2463,
// 16'h166e, 16'h0805, 16'hf96f, 16'heb20,
// 16'hdcfa, 16'hcfab, 16'hc357, 16'hb83d,
// 16'hae98, 16'ha69a, 16'ha06a, 16'h9c29,
// 16'h99f4, 16'h99c8, 16'h9bb5, 16'h9fa6,
// 16'ha58e, 16'had48, 16'hb6b4, 16'hc195,
// 16'hcdc2, 16'hdaec, 16'he8de, 16'hf740,
// 16'h05d6, 16'h144a, 16'h2256, 16'h2fb0,
// 16'h3c13, 16'h473b, 16'h50f8, 16'h5909,
// 16'h5f54, 16'h63aa, 16'h65ff, 16'h6640,
// 16'h6472, 16'h6097, 16'h5aca, 16'h5325,
// 16'h49cf, 16'h3efd, 16'h32e3, 16'h25bf,
// 16'h17db, 16'h0977, 16'hfae7, 16'hec6c,
// 16'hde5a, 16'hd0f7, 16'hc483, 16'hb94c,
// 16'haf7c, 16'ha751, 16'ha0f4, 16'h9c7f,
// 16'h9a14, 16'h99b5, 16'h9b6c, 16'h9f2a,
// 16'ha4e1, 16'hac6f, 16'hb5ae, 16'hc074,
// 16'hcc77, 16'hd998, 16'he76c, 16'hf5d1,
// 16'h045e, 16'h12de, 16'h20f3, 16'h2e66,
// 16'h3ae1, 16'h462f, 16'h5011, 16'h584e,
// 16'h5ec9, 16'h6352, 16'h65da, 16'h6654,
// 16'h64b5, 16'h6113, 16'h5b73, 16'h53fd,
// 16'h4ad0, 16'h4022, 16'h3425, 16'h2719,
// 16'h1947, 16'h0ae9, 16'hfc5e, 16'hedd8,
// 16'hdfbf, 16'hd240, 16'hc5ba, 16'hba57,
// 16'hb068, 16'ha80c, 16'ha182, 16'h9cdb,
// 16'h9a39, 16'h99a7, 16'h9b28, 16'h9eb4,
// 16'ha438, 16'hab9a, 16'hb4af, 16'hbf4f,
// 16'hcb3a, 16'hd839, 16'he607, 16'hf45a,
// 16'h02ec, 16'h116b, 16'h1f94, 16'h2d15,
// 16'h39af, 16'h451e, 16'h4f23, 16'h5793,
// 16'h5e36, 16'h62f5, 16'h65b3, 16'h665c,
// 16'h64fb, 16'h6183, 16'h5c1b, 16'h54d0,
// 16'h4bcd, 16'h4144, 16'h3564, 16'h2873,
// 16'h1aae, 16'h0c5f, 16'hfdcf, 16'hef4e,
// 16'he11c, 16'hd395, 16'hc6e9, 16'hbb6f,
// 16'hb152, 16'ha8d0, 16'ha213, 16'h9d3b,
// 16'h9a66, 16'h999c, 16'h9aeb, 16'h9e42,
// 16'ha394, 16'haaca, 16'hb3b3, 16'hbe2f,
// 16'hc9fc, 16'hd6e2, 16'he49e, 16'hf2e8,
// 16'h0175, 16'h0ffb, 16'h1e30, 16'h2bc5,
// 16'h3879, 16'h4408, 16'h4e34, 16'h56ce,
// 16'h5da2, 16'h6294, 16'h6581, 16'h6668,
// 16'h6530, 16'h61f8, 16'h5cb9, 16'h559f,
// 16'h4cc8, 16'h4260, 16'h36a3, 16'h29c9,
// 16'h1c15, 16'h0dd2, 16'hff44, 16'hf0be,
// 16'he283, 16'hd4e5, 16'hc822, 16'hbc84,
// 16'hb245, 16'ha995, 16'ha2aa, 16'h9da2,
// 16'h9a94, 16'h999b, 16'h9ab0, 16'h9dd5,
// 16'ha2f8, 16'ha9fa, 16'hb2bf, 16'hbd0f,
// 16'hc8c3, 16'hd58b, 16'he338, 16'hf176,
// 16'hfffe, 16'h0e8d, 16'h1cc7, 16'h2a74,
// 16'h373f, 16'h42f0, 16'h4d41, 16'h5605,
// 16'h5d0a, 16'h6229, 16'h6551, 16'h6665,
// 16'h656b, 16'h625f, 16'h5d57, 16'h5668,
// 16'h4dbd, 16'h437c, 16'h37dd, 16'h2b1c,
// 16'h1d7c, 16'h0f44, 16'h20b9, 16'hf232,
// 16'he3e5, 16'hd63d, 16'hc959, 16'hbda3,
// 16'hb336, 16'haa63, 16'ha343, 16'h9e0e,
// 16'h9aca, 16'h999c, 16'h9a7d, 16'h9d6d,
// 16'ha25e, 16'ha932, 16'hb1cb, 16'hbbf8,
// 16'hc788, 16'hd43a, 16'he1d2, 16'hf002,
// 16'hfe8e, 16'h0d14, 16'h1b67, 16'h291a,
// 16'h3606, 16'h41d1, 16'h4c4d, 16'h5535,
// 16'h5c6e, 16'h61bb, 16'h6519, 16'h6660,
// 16'h659e, 16'h62c0, 16'h5df3, 16'h572b,
// 16'h4eb1, 16'h448f, 16'h3918, 16'h2c6b,
// 16'h1ee4, 16'h10b2, 16'h0231, 16'hf3a1,
// 16'he552, 16'hd78d, 16'hca9d, 16'hbeba,
// 16'hb436, 16'hab2d, 16'ha3e8, 16'h9e79,
// 16'h9b09, 16'h99a1, 16'h9a50, 16'h9d09,
// 16'ha1ca, 16'ha86d, 16'hb0de, 16'hbae1,
// 16'hc652, 16'hd2ea, 16'he06d, 16'hee93,
// 16'hfd17, 16'h0ba3, 16'h19fc, 16'h27c4,
// 16'h34c8, 16'h40b0, 16'h4b51, 16'h5467,
// 16'h5bc7, 16'h614d, 16'h64d7, 16'h6659,
// 16'h65c8, 16'h6324, 16'h5e80, 16'h57f1,
// 16'h4f9b, 16'h45a6, 16'h3a49, 16'h2dbd,
// 16'h2044, 16'h1225, 16'h03a5, 16'hf514,
// 16'he6bb, 16'hd8e7, 16'hcbd9, 16'hbfe0,
// 16'hb52f, 16'hac03, 16'ha48e, 16'h9eec,
// 16'h9b4a, 16'h99ae, 16'h9a25, 16'h9caf,
// 16'ha136, 16'ha7b2, 16'hafee, 16'hb9d4,
// 16'hc51d, 16'hd19b, 16'hdf0c, 16'hed23,
// 16'hfba0, 16'h0a33, 16'h188f, 16'h266e,
// 16'h3383, 16'h3f90, 16'h4a4f, 16'h5395,
// 16'h5b1b, 16'h60da, 16'h6490, 16'h664d,
// 16'h65ed, 16'h637e, 16'h5f11, 16'h58a9,
// 16'h5089, 16'h46b1, 16'h3b7e, 16'h2f0a,
// 16'h21a4, 16'h1395, 16'h051a, 16'hf686,
// 16'he82a, 16'hda3b, 16'hcd23, 16'hc0fe,
// 16'hb635, 16'hacd8, 16'ha538, 16'h9f69,
// 16'h9b8c, 16'h99c3, 16'h99fe, 16'h9c57,
// 16'ha0ad, 16'ha6f5, 16'haf0a, 16'hb8c4,
// 16'hc3ec, 16'hd051, 16'hddaa, 16'hebb5,
// 16'hfa2c, 16'h08be, 16'h1723, 16'h2514,
// 16'h323e, 16'h3e6a, 16'h494e, 16'h52b6,
// 16'h5a74, 16'h6058, 16'h644d, 16'h6636,
// 16'h660d, 16'h63d8, 16'h5f93, 16'h596a,
// 16'h5165, 16'h47c5, 16'h3ca6, 16'h3059,
// 16'h2301, 16'h1506, 16'h068c, 16'hf7fe,
// 16'he991, 16'hdb9b, 16'hce65, 16'hc22b,
// 16'hb734, 16'hadb9, 16'ha5e4, 16'h9fe8,
// 16'h9bd9, 16'h99d7, 16'h99e1, 16'h9c03,
// 16'ha029, 16'ha63c, 16'hae2b, 16'hb7b5,
// 16'hc2c3, 16'hcf07, 16'hdc49, 16'hea4b,
// 16'hf8b3, 16'h074d, 16'h15b5, 16'h23b7,
// 16'h30f8, 16'h3d40, 16'h4847, 16'h51d8,
// 16'h59c2, 16'h5fd8, 16'h63fe, 16'h661e,
// 16'h6629, 16'h6427, 16'h6019, 16'h5a19,
// 16'h524b, 16'h48c9, 16'h3dd6, 16'h319c,
// 16'h2463, 16'h1670, 16'h0802, 16'hf973,
// 16'heafd, 16'hdcfa, 16'hcfac, 16'hc355,
// 16'hb840, 16'hae97, 16'ha69a, 16'ha068,
// 16'h9c2d, 16'h99ef, 16'h99ce, 16'h9baf,
// 16'h9fab, 16'ha58a, 16'had4c, 16'hb6b0,
// 16'hc198, 16'hcdbf, 16'hdaef, 16'he8db,
// 16'hf743, 16'h05d3, 16'h144d, 16'h2253,
// 16'h2fb3, 16'h3c10, 16'h473e, 16'h50f6,
// 16'h590b, 16'h5f52, 16'h63ac, 16'h65fe,
// 16'h6641, 16'h6470, 16'h609a, 16'h5ac7,
// 16'h5328, 16'h49cc, 16'h3eff, 16'h32e1,
// 16'h25c1, 16'h17da, 16'h0977, 16'hfae7,
// 16'hec6b, 16'hde5c, 16'hd0f4, 16'hc487,
// 16'hb948, 16'haf7e, 16'ha752, 16'ha0f1,
// 16'h9c83, 16'h9a0f, 16'h99b9, 16'h9b6a,
// 16'h9f2b, 16'ha4e2, 16'hac6c, 16'hb5b2,
// 16'hc06f, 16'hcc7d, 16'hd992, 16'he771,
// 16'hf5ce, 16'h0460, 16'h12db, 16'h20f6,
// 16'h2e64, 16'h3ae2, 16'h462f, 16'h500f,
// 16'h5851, 16'h5ec7, 16'h6352, 16'h65dc,
// 16'h6650, 16'h64bb, 16'h610d, 16'h5b78,
// 16'h53f9, 16'h4ad3, 16'h4020, 16'h3426,
// 16'h2719, 16'h1946, 16'h0aea, 16'hfc5d,
// 16'hedd9, 16'hdfbe, 16'hd240, 16'hc5ba,
// 16'hba58, 16'hb066, 16'ha80f, 16'ha17f,
// 16'h9cdc, 16'h9a39, 16'h99a8, 16'h9b27,
// 16'h9eb4, 16'ha439, 16'hab98, 16'hb4b2,
// 16'hbf4c, 16'hcb3c, 16'hd837, 16'he60a,
// 16'hf458, 16'h02ec, 16'h116b, 16'h1f94,
// 16'h2d15, 16'h39b1, 16'h451a, 16'h4f27,
// 16'h578f, 16'h5e39, 16'h62f4, 16'h65b3,
// 16'h665c, 16'h64fb, 16'h6182, 16'h5c1d,
// 16'h54cf, 16'h4bcd, 16'h4144, 16'h3563,
// 16'h2875, 16'h1aac, 16'h0c60, 16'hfdd0,
// 16'hef4b, 16'he120, 16'hd391, 16'hc6ec,
// 16'hbb6e, 16'hb151, 16'ha8d2, 16'ha211,
// 16'h9d3c, 16'h9a65, 16'h999e, 16'h9ae9,
// 16'h9e43, 16'ha394, 16'haac8, 16'hb3b7,
// 16'hbe2b, 16'hc9ff, 16'hd6e0, 16'he49e,
// 16'hf2e9, 16'h0174, 16'h0ffd, 16'h1e2e,
// 16'h2bc6, 16'h3878, 16'h4409, 16'h4e34,
// 16'h56ce, 16'h5da2, 16'h6293, 16'h6584,
// 16'h6663, 16'h6536, 16'h61f2, 16'h5cbe,
// 16'h559b, 16'h4ccc, 16'h425c, 16'h36a7,
// 16'h29c5, 16'h1c17, 16'h0dd2, 16'hff43,
// 16'hf0c1, 16'he27f, 16'hd4e8, 16'hc81f,
// 16'hbc87, 16'hb243, 16'ha996, 16'ha2aa,
// 16'h9da1, 16'h9a94, 16'h999d, 16'h9aae,
// 16'h9dd6, 16'ha2f7, 16'ha9fb, 16'hb2be,
// 16'hbd12, 16'hc8bf, 16'hd58e, 16'he337,
// 16'hf174, 16'h2003, 16'h0e87, 16'h1ccd,
// 16'h2a6f, 16'h3742, 16'h42ee, 16'h4d43,
// 16'h5603, 16'h5d0b, 16'h6229, 16'h6551,
// 16'h6665, 16'h656b, 16'h625e, 16'h5d58,
// 16'h5668, 16'h4dbd, 16'h437c, 16'h37dc,
// 16'h2b1e, 16'h1d7a, 16'h0f45, 16'h20b9,
// 16'hf230, 16'he3e9, 16'hd639, 16'hc95d,
// 16'hbd9e, 16'hb33b, 16'haa5e, 16'ha349,
// 16'h9e08, 16'h9acf, 16'h9998, 16'h9a7f,
// 16'h9d6d, 16'ha25e, 16'ha931, 16'hb1cd,
// 16'hbbf6, 16'hc789, 16'hd43a, 16'he1d1,
// 16'hf004, 16'hfe8c, 16'h0d17, 16'h1b63,
// 16'h291c, 16'h3606, 16'h41d1, 16'h4c4c,
// 16'h5537, 16'h5c6a, 16'h61c0, 16'h6515,
// 16'h6663, 16'h659b, 16'h62c3, 16'h5df0,
// 16'h572e, 16'h4eae, 16'h4493, 16'h3914,
// 16'h2c6e, 16'h1ee1, 16'h10b5, 16'h022e,
// 16'hf3a3, 16'he551, 16'hd78e, 16'hca9b,
// 16'hbebd, 16'hb431, 16'hab32, 16'ha3e5,
// 16'h9e7b, 16'h9b08, 16'h99a1, 16'h9a50,
// 16'h9d09, 16'ha1ca, 16'ha86e, 16'hb0dd,
// 16'hbae2, 16'hc651, 16'hd2ea, 16'he06d,
// 16'hee95, 16'hfd14, 16'h0ba6, 16'h19f8,
// 16'h27c9, 16'h34c3, 16'h40b5, 16'h4b4e,
// 16'h5467, 16'h5bc7, 16'h614e, 16'h64d5,
// 16'h665d, 16'h65c3, 16'h6327, 16'h5e7e,
// 16'h57f4, 16'h4f97, 16'h45aa, 16'h3a45,
// 16'h2dc1, 16'h2041, 16'h1228, 16'h03a2,
// 16'hf516, 16'he6bb, 16'hd8e5, 16'hcbdd,
// 16'hbfdd, 16'hb52f, 16'hac05, 16'ha48a,
// 16'h9ef1, 16'h9b47, 16'h99af, 16'h9a24,
// 16'h9caf, 16'ha137, 16'ha7b1, 16'hafef,
// 16'hb9d3, 16'hc51d, 16'hd19c, 16'hdf0a,
// 16'hed25, 16'hfba0, 16'h0a32, 16'h188f,
// 16'h266d, 16'h3385, 16'h3f8e, 16'h4a53,
// 16'h538f, 16'h5b21, 16'h60d3, 16'h6497,
// 16'h6648, 16'h65f0, 16'h637e, 16'h5f0d,
// 16'h58b0, 16'h5080, 16'h46bb, 16'h3b76,
// 16'h2f0d, 16'h21a5, 16'h1392, 16'h051e,
// 16'hf684, 16'he828, 16'hda3f, 16'hcd1d,
// 16'hc106, 16'hb62d, 16'hacdf, 16'ha533,
// 16'h9f6b, 16'h9b8d, 16'h99bf, 16'h9a03,
// 16'h9c54, 16'ha0ae, 16'ha6f5, 16'haf09,
// 16'hb8c4, 16'hc3ee, 16'hd04f, 16'hddab,
// 16'hebb4, 16'hfa2d, 16'h08bd, 16'h1725,
// 16'h2511, 16'h3242, 16'h3e66, 16'h4951,
// 16'h52b4, 16'h5a75, 16'h6059, 16'h644a,
// 16'h6639, 16'h660c, 16'h63d7, 16'h5f96,
// 16'h5965, 16'h5169, 16'h47c3, 16'h3ca8,
// 16'h3057, 16'h2303, 16'h1504, 16'h068d,
// 16'hf7ff, 16'he98e, 16'hdba0, 16'hce5f,
// 16'hc230, 16'hb732, 16'hadb9, 16'ha5e5,
// 16'h9fe6, 16'h9bdb, 16'h99d7, 16'h99e0,
// 16'h9c05, 16'ha025, 16'ha641, 16'hae27,
// 16'hb7b7, 16'hc2c4, 16'hcf03, 16'hdc4f,
// 16'hea45, 16'hf8b8, 16'h0749, 16'h15b8,
// 16'h23b5, 16'h30fa, 16'h3d3e, 16'h4848,
// 16'h51d9, 16'h59bf, 16'h5fdc, 16'h63fa,
// 16'h6620, 16'h662a, 16'h6424, 16'h601c,
// 16'h5a18, 16'h5249, 16'h48cc, 16'h3dd3,
// 16'h319f, 16'h2461, 16'h1671, 16'h0801,
// 16'hf973, 16'heafe, 16'hdcfa, 16'hcfac,
// 16'hc356, 16'hb83e, 16'hae97, 16'ha69b,
// 16'ha069, 16'h9c2c, 16'h99f0, 16'h99cb,
// 16'h9bb2, 16'h9fa9, 16'ha58c, 16'had4a,
// 16'hb6b2, 16'hc196, 16'hcdc2, 16'hdaec,
// 16'he8dd, 16'hf742, 16'h05d4, 16'h144c,
// 16'h2254, 16'h2fb3, 16'h3c0f, 16'h473f,
// 16'h50f5, 16'h590a, 16'h5f56, 16'h63a7,
// 16'h6602, 16'h663e, 16'h6473, 16'h6096,
// 16'h5acc, 16'h5323, 16'h49d0, 16'h3efe,
// 16'h32e0, 16'h25c2, 16'h17d9, 16'h0978,
// 16'hfae6, 16'hec6d, 16'hde59, 16'hd0f8,
// 16'hc482, 16'hb94d, 16'haf79, 16'ha756,
// 16'ha0ef, 16'h9c84, 16'h9a0f, 16'h99b8,
// 16'h9b6b, 16'h9f2a, 16'ha4e2, 16'hac6e,
// 16'hb5af, 16'hc071, 16'hcc7c, 16'hd992,
// 16'he772, 16'hf5cc, 16'h0461, 16'h12dc,
// 16'h20f4, 16'h2e66, 16'h3ae1, 16'h462e,
// 16'h5012, 16'h584d, 16'h5eca, 16'h6351,
// 16'h65dc, 16'h6651, 16'h64b9, 16'h610f,
// 16'h5b76, 16'h53fa, 16'h4ad4, 16'h401e,
// 16'h3428, 16'h2717, 16'h1947, 16'h0aeb,
// 16'hfc5b, 16'heddb, 16'hdfbd, 16'hd240,
// 16'hc5ba, 16'hba58, 16'hb066, 16'ha810,
// 16'ha17e, 16'h9cdc, 16'h9a39, 16'h99a8,
// 16'h9b27, 16'h9eb4, 16'ha439, 16'hab98,
// 16'hb4b2, 16'hbf4c, 16'hcb3b, 16'hd839,
// 16'he608, 16'hf459, 16'h02ec, 16'h116b,
// 16'h1f94, 16'h2d15, 16'h39b0, 16'h451c,
// 16'h4f25, 16'h5790, 16'h5e39, 16'h62f4,
// 16'h65b2, 16'h665f, 16'h64f6, 16'h6187,
// 16'h5c1a, 16'h54ce, 16'h4bd1, 16'h413f,
// 16'h3569, 16'h286f, 16'h1ab0, 16'h0c5e,
// 16'hfdd0, 16'hef4c, 16'he11f, 16'hd392,
// 16'hc6ec, 16'hbb6c, 16'hb154, 16'ha8d0,
// 16'ha212, 16'h9d3c, 16'h9a64, 16'h999f,
// 16'h9ae8, 16'h9e44, 16'ha393, 16'haaca,
// 16'hb3b4, 16'hbe2d, 16'hc9fe, 16'hd6e0,
// 16'he4a0, 16'hf2e6, 16'h0176, 16'h0ffd,
// 16'h1e2d, 16'h2bc7, 16'h3878, 16'h4407,
// 16'h4e38, 16'h56c9, 16'h5da7, 16'h628f,
// 16'h6586, 16'h6663, 16'h6534, 16'h61f5,
// 16'h5cbb, 16'h559f, 16'h4cc7, 16'h4260,
// 16'h36a4, 16'h29c7, 16'h1c16, 16'h0dd3,
// 16'hff42, 16'hf0c1, 16'he27f, 16'hd4e9,
// 16'hc81e, 16'hbc89, 16'hb240, 16'ha998,
// 16'ha2a9, 16'h9da1, 16'h9a96, 16'h999b,
// 16'h9aaf, 16'h9dd5, 16'ha2f8, 16'ha9fa,
// 16'hb2c0, 16'hbd0f, 16'hc8c2, 16'hd58b,
// 16'he33a, 16'hf172, 16'h2003, 16'h0e89,
// 16'h1cc8, 16'h2a76, 16'h373c, 16'h42f2,
// 16'h4d40, 16'h5606, 16'h5d08, 16'h622d,
// 16'h654d, 16'h6668, 16'h6569, 16'h625f,
// 16'h5d58, 16'h5668, 16'h4dbe, 16'h4379,
// 16'h37e0, 16'h2b1a, 16'h1d7d, 16'h0f43,
// 16'h20ba, 16'hf230, 16'he3e9, 16'hd639,
// 16'hc95c, 16'hbda0, 16'hb339, 16'haa60,
// 16'ha347, 16'h9e0a, 16'h9acc, 16'h999c,
// 16'h9a7d, 16'h9d6c, 16'ha260, 16'ha930,
// 16'hb1cc, 16'hbbf8, 16'hc788, 16'hd43a,
// 16'he1d1, 16'hf005, 16'hfe89, 16'h0d1a,
// 16'h1b62, 16'h291d, 16'h3604, 16'h41d2,
// 16'h4c4b, 16'h553a, 16'h5c68, 16'h61c1,
// 16'h6513, 16'h6665, 16'h6599, 16'h62c6,
// 16'h5dee, 16'h572e, 16'h4eaf, 16'h4492,
// 16'h3914, 16'h2c6f, 16'h1ee0, 16'h10b5,
// 16'h0230, 16'hf3a1, 16'he552, 16'hd78d,
// 16'hca9c, 16'hbebd, 16'hb431, 16'hab32,
// 16'ha3e4, 16'h9e7c, 16'h9b07, 16'h99a3,
// 16'h9a4c, 16'h9d0e, 16'ha1c5, 16'ha873,
// 16'hb0d8, 16'hbae5, 16'hc650, 16'hd2ea,
// 16'he06e, 16'hee94, 16'hfd13, 16'h0ba9,
// 16'h19f5, 16'h27cb, 16'h34c2, 16'h40b4,
// 16'h4b50, 16'h5466, 16'h5bc8, 16'h614c,
// 16'h64d8, 16'h6659, 16'h65c7, 16'h6324,
// 16'h5e81, 16'h57f1, 16'h4f9a, 16'h45a6,
// 16'h3a4a, 16'h2dbd, 16'h2045, 16'h1222,
// 16'h03a8, 16'hf511, 16'he6c0, 16'hd8e1,
// 16'hcbdf, 16'hbfdc, 16'hb530, 16'hac04,
// 16'ha48b, 16'h9ef0, 16'h9b48, 16'h99ae,
// 16'h9a25, 16'h9cad, 16'ha13a, 16'ha7ad,
// 16'haff5, 16'hb9cd, 16'hc521, 16'hd19a,
// 16'hdf0b, 16'hed25, 16'hfba0, 16'h0a31,
// 16'h1892, 16'h2669, 16'h3388, 16'h3f8d,
// 16'h4a52, 16'h5391, 16'h5b1e, 16'h60d7,
// 16'h6494, 16'h664b, 16'h65eb, 16'h6383,
// 16'h5f0a, 16'h58b2, 16'h5080, 16'h46b8,
// 16'h3b7a, 16'h2f0b, 16'h21a4, 16'h1396,
// 16'h0518, 16'hf68a, 16'he825, 16'hda3f,
// 16'hcd1f, 16'hc103, 16'hb630, 16'hacdc,
// 16'ha535, 16'h9f69, 16'h9b90, 16'h99bd,
// 16'h9a03, 16'h9c54, 16'ha0ae, 16'ha6f5,
// 16'haf0a, 16'hb8c3, 16'hc3ee, 16'hd050,
// 16'hddaa, 16'hebb5, 16'hfa2c, 16'h08bc,
// 16'h1728, 16'h250e, 16'h3243, 16'h3e67,
// 16'h494e, 16'h52b9, 16'h5a70, 16'h605c,
// 16'h6448, 16'h663b, 16'h660a, 16'h63da,
// 16'h5f91, 16'h596a, 16'h5166, 16'h47c4,
// 16'h3ca8, 16'h3055, 16'h2305, 16'h1503,
// 16'h068f, 16'hf7fb, 16'he994, 16'hdb98,
// 16'hce69, 16'hc225, 16'hb73b, 16'hadb3,
// 16'ha5e9, 16'h9fe4, 16'h9bdb, 16'h99d6,
// 16'h99e2, 16'h9c04, 16'ha025, 16'ha640,
// 16'hae27, 16'hb7b9, 16'hc2c1, 16'hcf07,
// 16'hdc4a, 16'hea48, 16'hf8b7, 16'h0749,
// 16'h15b9, 16'h23b5, 16'h30f7, 16'h3d43,
// 16'h4843, 16'h51dc, 16'h59bf, 16'h5fda,
// 16'h63fd, 16'h661e, 16'h6629, 16'h6427,
// 16'h6018, 16'h5a1c, 16'h5247, 16'h48cc,
// 16'h3dd4, 16'h319d, 16'h2463, 16'h166f,
// 16'h0804, 16'hf970, 16'heb20, 16'hdcf8,
// 16'hcfad, 16'hc356, 16'hb83e, 16'hae98,
// 16'ha699, 16'ha06a, 16'h9c2b, 16'h99f1,
// 16'h99ca, 16'h9bb4, 16'h9fa6, 16'ha58e,
// 16'had48, 16'hb6b3, 16'hc196, 16'hcdc1,
// 16'hdaed, 16'he8dd, 16'hf740, 16'h05d7,
// 16'h1449, 16'h2257, 16'h2faf, 16'h3c12,
// 16'h473e, 16'h50f5, 16'h590c, 16'h5f51,
// 16'h63ac, 16'h65fe, 16'h6641, 16'h6471,
// 16'h6097, 16'h5acc, 16'h5322, 16'h49d2,
// 16'h3efa, 16'h32e4, 16'h25c0, 16'h17d9,
// 16'h0979, 16'hfae5, 16'hec6d, 16'hde5a,
// 16'hd0f6, 16'hc485, 16'hb94a, 16'haf7c,
// 16'ha753, 16'ha0f1, 16'h9c83, 16'h9a10,
// 16'h99b7, 16'h9b6b, 16'h9f2b, 16'ha4e0,
// 16'hac70, 16'hb5ad, 16'hc073, 16'hcc7a,
// 16'hd995, 16'he76e, 16'hf5d0, 16'h045e,
// 16'h12dc, 16'h20f8, 16'h2e60, 16'h3ae7,
// 16'h462a, 16'h5012, 16'h5850, 16'h5ec6,
// 16'h6356, 16'h65d6, 16'h6656, 16'h64b4,
// 16'h6114, 16'h5b73, 16'h53fd, 16'h4acf,
// 16'h4023, 16'h3423, 16'h271e, 16'h1940,
// 16'h0af1, 16'hfc55, 16'hede1, 16'hdfb8,
// 16'hd244, 16'hc5b7, 16'hba5a, 16'hb065,
// 16'ha810, 16'ha17e, 16'h9cdc, 16'h9a3a,
// 16'h99a6, 16'h9b2a, 16'h9eb1, 16'ha43b,
// 16'hab98, 16'hb4b0, 16'hbf4f, 16'hcb39,
// 16'hd83a, 16'he608, 16'hf458, 16'h02ed,
// 16'h116b, 16'h1f93, 16'h2d16, 16'h39b0,
// 16'h451b, 16'h4f27, 16'h578e, 16'h5e3a,
// 16'h62f4, 16'h65b1, 16'h6660, 16'h64f6,
// 16'h6187, 16'h5c1a, 16'h54ce, 16'h4bd0,
// 16'h4141, 16'h3567, 16'h2871, 16'h1aaf,
// 16'h0c5e, 16'hfdd1, 16'hef4b, 16'he120,
// 16'hd390, 16'hc6ed, 16'hbb6e, 16'hb151,
// 16'ha8d2, 16'ha211, 16'h9d3b, 16'h9a67,
// 16'h999c, 16'h9aeb, 16'h9e41, 16'ha395,
// 16'haaca, 16'hb3b2, 16'hbe31, 16'hc9f9,
// 16'hd6e5, 16'he49c, 16'hf2e9, 16'h0174,
// 16'h0ffd, 16'h1e2f, 16'h2bc4, 16'h387c,
// 16'h4404, 16'h4e38, 16'h56cc, 16'h5da2,
// 16'h6295, 16'h6580, 16'h6668, 16'h6531,
// 16'h61f7, 16'h5cb9, 16'h55a1, 16'h4cc5,
// 16'h4263, 16'h369f, 16'h29cd, 16'h1c12,
// 16'h0dd4, 16'hff44, 16'hf0bc, 16'he286,
// 16'hd4e2, 16'hc824, 16'hbc84, 16'hb244,
// 16'ha996, 16'ha2ab, 16'h9d9e, 16'h9a99,
// 16'h9997, 16'h9ab4, 16'h9dd2, 16'ha2f9,
// 16'ha9fa, 16'hb2bd, 16'hbd14, 16'hc8bd,
// 16'hd590, 16'he335, 16'hf176, 16'h2001,
// 16'h0e89, 16'h1cca, 16'h2a72, 16'h3740,
// 16'h42f0, 16'h4d40, 16'h5607, 16'h5d07,
// 16'h622d, 16'h654e, 16'h6667, 16'h6569,
// 16'h6260, 16'h5d57, 16'h5669, 16'h4dbd,
// 16'h437a, 16'h37df, 16'h2b1a, 16'h1d7e,
// 16'h0f43, 16'h20b9, 16'hf231, 16'he3e9,
// 16'hd637, 16'hc960, 16'hbd9c, 16'hb33a,
// 16'haa63, 16'ha342, 16'h9e0f, 16'h9ac9,
// 16'h999d, 16'h9a7b, 16'h9d70, 16'ha25b,
// 16'ha934, 16'hb1cb, 16'hbbf6, 16'hc78a,
// 16'hd438, 16'he1d4, 16'hf002, 16'hfe8b,
// 16'h0d18, 16'h1b62, 16'h291f, 16'h3603,
// 16'h41d3, 16'h4c49, 16'h553a, 16'h5c69,
// 16'h61c1, 16'h6513, 16'h6666, 16'h6596,
// 16'h62c9, 16'h5deb, 16'h5732, 16'h4eab,
// 16'h4495, 16'h3912, 16'h2c70, 16'h1ee0,
// 16'h10b4, 16'h0231, 16'hf3a0, 16'he553,
// 16'hd78e, 16'hca99, 16'hbec0, 16'hb42f,
// 16'hab33, 16'ha3e4, 16'h9e7c, 16'h9b07,
// 16'h99a2, 16'h9a4e, 16'h9d0c, 16'ha1c7,
// 16'ha871, 16'hb0d9, 16'hbae5, 16'hc650,
// 16'hd2eb, 16'he06c, 16'hee94, 16'hfd16,
// 16'h0ba4, 16'h19fb, 16'h27c5, 16'h34c7,
// 16'h40b1, 16'h4b51, 16'h5466, 16'h5bc7,
// 16'h614e, 16'h64d6, 16'h665b, 16'h65c4,
// 16'h6327, 16'h5e7e, 16'h57f3, 16'h4f9a,
// 16'h45a5, 16'h3a4a, 16'h2dbd, 16'h2044,
// 16'h1225, 16'h03a4, 16'hf516, 16'he6ba,
// 16'hd8e7, 16'hcbd9, 16'hbfe1, 16'hb52d,
// 16'hac06, 16'ha48a, 16'h9ef0, 16'h9b48,
// 16'h99af, 16'h9a24, 16'h9cae, 16'ha139,
// 16'ha7af, 16'haff1, 16'hb9d1, 16'hc51e,
// 16'hd19d, 16'hdf09, 16'hed25, 16'hfba0,
// 16'h0a31, 16'h1893, 16'h2668, 16'h3389,
// 16'h3f8b, 16'h4a55, 16'h538e, 16'h5b21,
// 16'h60d5, 16'h6494, 16'h664c, 16'h65eb,
// 16'h6382, 16'h5f0b, 16'h58b1, 16'h5081,
// 16'h46b8, 16'h3b79, 16'h2f0b, 16'h21a6,
// 16'h1393, 16'h051b, 16'hf688, 16'he825,
// 16'hda40, 16'hcd1e, 16'hc105, 16'hb62e,
// 16'hacde, 16'ha533, 16'h9f6a, 16'h9b90,
// 16'h99bd, 16'h9a03, 16'h9c54, 16'ha0ae,
// 16'ha6f6, 16'haf09, 16'hb8c2, 16'hc3f1,
// 16'hd04c, 16'hddae, 16'hebb2, 16'hfa2d,
// 16'h08be, 16'h1723, 16'h2514, 16'h323d,
// 16'h3e6b, 16'h494e, 16'h52b5, 16'h5a75,
// 16'h6057, 16'h644d, 16'h6637, 16'h660e,
// 16'h63d5, 16'h5f96, 16'h5966, 16'h5169,
// 16'h47c2, 16'h3ca9, 16'h3056, 16'h2304,
// 16'h1502, 16'h068f, 16'hf7fd, 16'he990,
// 16'hdb9f, 16'hce60, 16'hc22d, 16'hb735,
// 16'hadb7, 16'ha5e6, 16'h9fe7, 16'h9bd9,
// 16'h99d6, 16'h99e3, 16'h9c02, 16'ha027,
// 16'ha640, 16'hae26, 16'hb7b9, 16'hc2c1,
// 16'hcf07, 16'hdc4a, 16'hea4b, 16'hf8b2,
// 16'h074e, 16'h15b4, 16'h23b8, 16'h30f8,
// 16'h3d40, 16'h4846, 16'h51da, 16'h59bf,
// 16'h5fdc, 16'h63fa, 16'h6621, 16'h6626,
// 16'h6429, 16'h6018, 16'h5a1b, 16'h5248,
// 16'h48cb, 16'h3dd4, 16'h319e, 16'h2463,
// 16'h166e, 16'h0805, 16'hf96f, 16'heb01,
// 16'hdcf9, 16'hcfab, 16'hc357, 16'hb83e,
// 16'hae97, 16'ha69b, 16'ha068, 16'h9c2d,
// 16'h99f0, 16'h99cb, 16'h9bb2, 16'h9fa8,
// 16'ha58d, 16'had49, 16'hb6b3, 16'hc195,
// 16'hcdc2, 16'hdaec, 16'he8de, 16'hf740,
// 16'h05d6, 16'h144b, 16'h2254, 16'h2fb3,
// 16'h3c0f, 16'h473f, 16'h50f7, 16'h5908,
// 16'h5f56, 16'h63a6, 16'h6604, 16'h663d,
// 16'h6474, 16'h6096, 16'h5ac9, 16'h5327,
// 16'h49cd, 16'h3f20, 16'h32df, 16'h25c3,
// 16'h17d6, 16'h097d, 16'hfae1, 16'hec70,
// 16'hde59, 16'hd0f4, 16'hc488, 16'hb948,
// 16'haf7d, 16'ha752, 16'ha0f2, 16'h9c81,
// 16'h9a12, 16'h99b7, 16'h9b6a, 16'h9f2c,
// 16'ha4df, 16'hac70, 16'hb5af, 16'hc072,
// 16'hcc7a, 16'hd994, 16'he770, 16'hf5ce,
// 16'h0461, 16'h12da, 16'h20f7, 16'h2e63,
// 16'h3ae4, 16'h462c, 16'h5012, 16'h584d,
// 16'h5ecc, 16'h634e, 16'h65de, 16'h6650,
// 16'h64b8, 16'h6111, 16'h5b75, 16'h53fb,
// 16'h4ad2, 16'h4020, 16'h3426, 16'h271a,
// 16'h1945, 16'h0aec, 16'hfc59, 16'hedde,
// 16'hdfb9, 16'hd246, 16'hc5b5, 16'hba5a,
// 16'hb065, 16'ha810, 16'ha17e, 16'h9cdf,
// 16'h9a35, 16'h99ab, 16'h9b24, 16'h9eb7,
// 16'ha437, 16'hab9a, 16'hb4b0, 16'hbf4d,
// 16'hcb3b, 16'hd839, 16'he607, 16'hf45a,
// 16'h02ec, 16'h116b, 16'h1f93, 16'h2d16,
// 16'h39af, 16'h451d, 16'h4f25, 16'h5790,
// 16'h5e38, 16'h62f6, 16'h65af, 16'h6662,
// 16'h64f3, 16'h618c, 16'h5c13, 16'h54d6,
// 16'h4bc9, 16'h4146, 16'h3563, 16'h2874,
// 16'h1aad, 16'h0c5f, 16'hfdd1, 16'hef4a,
// 16'he121, 16'hd390, 16'hc6ee, 16'hbb6b,
// 16'hb154, 16'ha8d0, 16'ha212, 16'h9d3c,
// 16'h9a65, 16'h999d, 16'h9aea, 16'h9e43,
// 16'ha394, 16'haac9, 16'hb3b4, 16'hbe2e,
// 16'hc9fc, 16'hd6e3, 16'he49d, 16'hf2e9,
// 16'h0174, 16'h0ffc, 16'h1e2f, 16'h2bc5,
// 16'h387a, 16'h4407, 16'h4e36, 16'h56cb,
// 16'h5da5, 16'h6290, 16'h6587, 16'h6661,
// 16'h6536, 16'h61f4, 16'h5cba, 16'h55a1,
// 16'h4cc5, 16'h4262, 16'h36a2, 16'h29c8,
// 16'h1c17, 16'h0dd0, 16'hff46, 16'hf0bd,
// 16'he283, 16'hd4e5, 16'hc822, 16'hbc84,
// 16'hb246, 16'ha994, 16'ha2ab, 16'h9da0,
// 16'h9a95, 16'h999c, 16'h9aaf, 16'h9dd6,
// 16'ha2f6, 16'ha9fb, 16'hb2bf, 16'hbd10,
// 16'hc8c1, 16'hd58d, 16'he336, 16'hf177,
// 16'hfffe, 16'h0e8d, 16'h1cc7, 16'h2a73,
// 16'h3740, 16'h42ef, 16'h4d42, 16'h5605,
// 16'h5d09, 16'h622b, 16'h654f, 16'h6666,
// 16'h656b, 16'h625e, 16'h5d59, 16'h5667,
// 16'h4dbe, 16'h437a, 16'h37de, 16'h2b1c,
// 16'h1d7c, 16'h0f43, 16'h20bb, 16'hf22e,
// 16'he3eb, 16'hd638, 16'hc95c, 16'hbda1,
// 16'hb336, 16'haa64, 16'ha344, 16'h9e0c,
// 16'h9acb, 16'h999c, 16'h9a7c, 16'h9d6f,
// 16'ha25c, 16'ha933, 16'hb1ca, 16'hbbfa,
// 16'hc786, 16'hd43b, 16'he1d1, 16'hf004,
// 16'hfe8b, 16'h0d19, 16'h1b60, 16'h2920,
// 16'h3602, 16'h41d5, 16'h4c47, 16'h553d,
// 16'h5c66, 16'h61c1, 16'h6516, 16'h6660,
// 16'h659e, 16'h62c2, 16'h5df0, 16'h572e,
// 16'h4eaf, 16'h4490, 16'h3917, 16'h2c6c,
// 16'h1ee3, 16'h10b2, 16'h0232, 16'hf39f,
// 16'he554, 16'hd78c, 16'hca9c, 16'hbebc,
// 16'hb433, 16'hab30, 16'ha3e6, 16'h9e7b,
// 16'h9b07, 16'h99a3, 16'h9a4e, 16'h9d0b,
// 16'ha1c8, 16'ha870, 16'hb0da, 16'hbae5,
// 16'hc650, 16'hd2ea, 16'he06e, 16'hee92,
// 16'hfd16, 16'h0ba6, 16'h19f9, 16'h27c7,
// 16'h34c5, 16'h40b3, 16'h4b4f, 16'h5467,
// 16'h5bc8, 16'h614c, 16'h64d8, 16'h6659,
// 16'h65c6, 16'h6325, 16'h5e81, 16'h57ef,
// 16'h4f9e, 16'h45a1, 16'h3a4e, 16'h2dba,
// 16'h2047, 16'h1223, 16'h03a4, 16'hf517,
// 16'he6b9, 16'hd8e8, 16'hcbd9, 16'hbfdf,
// 16'hb530, 16'hac04, 16'ha48b, 16'h9eef,
// 16'h9b48, 16'h99af, 16'h9a25, 16'h9cae,
// 16'ha138, 16'ha7af, 16'haff2, 16'hb9d0,
// 16'hc520, 16'hd199, 16'hdf0d, 16'hed22,
// 16'hfba2, 16'h0a31, 16'h188f, 16'h266f,
// 16'h3382, 16'h3f91, 16'h4a4f, 16'h5393,
// 16'h5b1e, 16'h60d6, 16'h6495, 16'h664a,
// 16'h65ec, 16'h6382, 16'h5f0b, 16'h58b0,
// 16'h5083, 16'h46b5, 16'h3b7c, 16'h2f09,
// 16'h21a7, 16'h1393, 16'h051a, 16'hf688,
// 16'he826, 16'hda3f, 16'hcd20, 16'hc101,
// 16'hb632, 16'hacda, 16'ha537, 16'h9f68,
// 16'h9b8f, 16'h99c0, 16'h9a01, 16'h9c54,
// 16'ha0ae, 16'ha6f5, 16'haf0b, 16'hb8c2,
// 16'hc3ef, 16'hd04e, 16'hddac, 16'hebb4,
// 16'hfa2c, 16'h08bd, 16'h1726, 16'h2511,
// 16'h3240, 16'h3e69, 16'h494d, 16'h52b9,
// 16'h5a70, 16'h605d, 16'h6448, 16'h6639,
// 16'h660e, 16'h63d4, 16'h5f99, 16'h5963,
// 16'h516a, 16'h47c2, 16'h3ca9, 16'h3057,
// 16'h2301, 16'h1506, 16'h068b, 16'hf801,
// 16'he98e, 16'hdb9e, 16'hce62, 16'hc22c,
// 16'hb735, 16'hadb8, 16'ha5e5, 16'h9fe7,
// 16'h9bda, 16'h99d6, 16'h99e2, 16'h9c03,
// 16'ha028, 16'ha63e, 16'hae28, 16'hb7b8,
// 16'hc2c1, 16'hcf08, 16'hdc4a, 16'hea48,
// 16'hf8b7, 16'h0749, 16'h15b8, 16'h23b5,
// 16'h30f9, 16'h3d40, 16'h4847, 16'h51d8,
// 16'h59c2, 16'h5fd6, 16'h6402, 16'h661a,
// 16'h662d, 16'h6423, 16'h601b, 16'h5a1a,
// 16'h5249, 16'h48ca, 16'h3dd6, 16'h319b,
// 16'h2465, 16'h166e, 16'h0804, 16'hf970,
// 16'heb20, 16'hdcf8, 16'hcfad, 16'hc356,
// 16'hb83d, 16'hae9a, 16'ha696, 16'ha06e,
// 16'h9c27, 16'h99f5, 16'h99c8, 16'h9bb4,
// 16'h9fa7, 16'ha58d, 16'had49, 16'hb6b3,
// 16'hc197, 16'hcdbf, 16'hdaef, 16'he8db,
// 16'hf742, 16'h05d6, 16'h1449, 16'h2257,
// 16'h2fb0, 16'h3c12, 16'h473d, 16'h50f6,
// 16'h590b, 16'h5f52, 16'h63ac, 16'h65fe,
// 16'h6640, 16'h6473, 16'h6096, 16'h5aca,
// 16'h5326, 16'h49ce, 16'h3efe, 16'h32e1,
// 16'h25c0, 16'h17db, 16'h0978, 16'hfae5,
// 16'hec6c, 16'hde5c, 16'hd0f4, 16'hc487,
// 16'hb948, 16'haf7d, 16'ha754, 16'ha0ef,
// 16'h9c84, 16'h9a0f, 16'h99b9, 16'h9b6a,
// 16'h9f2a, 16'ha4e2, 16'hac6d, 16'hb5b1,
// 16'hc070, 16'hcc7c, 16'hd993, 16'he770,
// 16'hf5ce, 16'h0461, 16'h12da, 16'h20f7,
// 16'h2e63, 16'h3ae2, 16'h4631, 16'h500c,
// 16'h5853, 16'h5ec6, 16'h6352, 16'h65dd,
// 16'h664f, 16'h64bb, 16'h610d, 16'h5b78,
// 16'h53fa, 16'h4ad2, 16'h4021, 16'h3424,
// 16'h271c, 16'h1944, 16'h0aec, 16'hfc5a,
// 16'heddc, 16'hdfbc, 16'hd243, 16'hc5b7,
// 16'hba58, 16'hb068, 16'ha80c, 16'ha183,
// 16'h9cd9, 16'h9a3a, 16'h99a8, 16'h9b25,
// 16'h9eb7, 16'ha436, 16'hab9b, 16'hb4af,
// 16'hbf4e, 16'hcb3a, 16'hd83a, 16'he607,
// 16'hf459, 16'h02ed, 16'h116a, 16'h1f95,
// 16'h2d15, 16'h39af, 16'h451d, 16'h4f26,
// 16'h578e, 16'h5e3b, 16'h62f3, 16'h65b1,
// 16'h6661, 16'h64f4, 16'h618a, 16'h5c16,
// 16'h54d2, 16'h4bcd, 16'h4142, 16'h3567,
// 16'h2870, 16'h1ab1, 16'h0c5c, 16'hfdd2,
// 16'hef4b, 16'he11f, 16'hd393, 16'hc6ea,
// 16'hbb6e, 16'hb153, 16'ha8d0, 16'ha213,
// 16'h9d3a, 16'h9a66, 16'h999d, 16'h9ae9,
// 16'h9e45, 16'ha391, 16'haacc, 16'hb3b2,
// 16'hbe30, 16'hc9f9, 16'hd6e6, 16'he49a,
// 16'hf2ec, 16'h0173, 16'h0ffc, 16'h1e2f,
// 16'h2bc5, 16'h387a, 16'h4408, 16'h4e34,
// 16'h56ce, 16'h5da2, 16'h6294, 16'h6582,
// 16'h6665, 16'h6534, 16'h61f5, 16'h5cbb,
// 16'h559f, 16'h4cc6, 16'h4261, 16'h36a4,
// 16'h29c6, 16'h1c19, 16'h0dce, 16'hff47,
// 16'hf0bc, 16'he284, 16'hd4e4, 16'hc822,
// 16'hbc86, 16'hb241, 16'ha99a, 16'ha2a6,
// 16'h9da3, 16'h9a95, 16'h9999, 16'h9ab2,
// 16'h9dd5, 16'ha2f6, 16'ha9fc, 16'hb2bd,
// 16'hbd12, 16'hc8c0, 16'hd58d, 16'he337,
// 16'hf175, 16'h2001, 16'h0e8a, 16'h1cc8,
// 16'h2a76, 16'h373b, 16'h42f3, 16'h4d3f,
// 16'h5608, 16'h5d06, 16'h622e, 16'h654c,
// 16'h6669, 16'h6569, 16'h6260, 16'h5d55,
// 16'h566b, 16'h4dbb, 16'h437d, 16'h37dd,
// 16'h2b1b, 16'h1d7d, 16'h0f43, 16'h20ba,
// 16'hf231, 16'he3e7, 16'hd63a, 16'hc95d,
// 16'hbd9e, 16'hb33b, 16'haa5e, 16'ha349,
// 16'h9e07, 16'h9ad1, 16'h9997, 16'h9a7f,
// 16'h9d6d, 16'ha25d, 16'ha933, 16'hb1cb,
// 16'hbbf8, 16'hc787, 16'hd43b, 16'he1d1,
// 16'hf004, 16'hfe8b, 16'h0d18, 16'h1b62,
// 16'h291e, 16'h3604, 16'h41d2, 16'h4c4b,
// 16'h5538, 16'h5c6a, 16'h61c0, 16'h6515,
// 16'h6662, 16'h659b, 16'h62c5, 16'h5dee,
// 16'h572f, 16'h4ead, 16'h4493, 16'h3915,
// 16'h2c6e, 16'h1ee0, 16'h10b5, 16'h022f,
// 16'hf3a3, 16'he550, 16'hd78f, 16'hca9a,
// 16'hbebe, 16'hb431, 16'hab32, 16'ha3e4,
// 16'h9e7c, 16'h9b07, 16'h99a2, 16'h9a4f,
// 16'h9d0b, 16'ha1c7, 16'ha871, 16'hb0d9,
// 16'hbae6, 16'hc64f, 16'hd2eb, 16'he06c,
// 16'hee95, 16'hfd14, 16'h0ba7, 16'h19f7,
// 16'h27c9, 16'h34c3, 16'h40b5, 16'h4b4e,
// 16'h5468, 16'h5bc6, 16'h614d, 16'h64d9,
// 16'h6657, 16'h65c9, 16'h6323, 16'h5e80,
// 16'h57f3, 16'h4f98, 16'h45a8, 16'h3a48,
// 16'h2dbe, 16'h2044, 16'h1224, 16'h03a6,
// 16'hf513, 16'he6bd, 16'hd8e5, 16'hcbda,
// 16'hbfe0, 16'hb52f, 16'hac02, 16'ha490,
// 16'h9ee9, 16'h9b4d, 16'h99ac, 16'h9a26,
// 16'h9cad, 16'ha139, 16'ha7af, 16'haff1,
// 16'hb9d1, 16'hc51f, 16'hd19a, 16'hdf0c,
// 16'hed24, 16'hfb9f, 16'h0a33, 16'h1890,
// 16'h266c, 16'h3385, 16'h3f8f, 16'h4a51,
// 16'h5391, 16'h5b20, 16'h60d3, 16'h6498,
// 16'h6647, 16'h65f1, 16'h637b, 16'h5f12,
// 16'h58ab, 16'h5084, 16'h46b8, 16'h3b77,
// 16'h2f0e, 16'h21a4, 16'h1394, 16'h051a,
// 16'hf688, 16'he825, 16'hda42, 16'hcd1c,
// 16'hc105, 16'hb62e, 16'hacdd, 16'ha535,
// 16'h9f6a, 16'h9b8d, 16'h99c1, 16'h99ff,
// 16'h9c58, 16'ha0aa, 16'ha6f9, 16'haf06,
// 16'hb8c7, 16'hc3ea, 16'hd053, 16'hdda8,
// 16'hebb7, 16'hfa2a, 16'h08be, 16'h1725,
// 16'h2512, 16'h323f, 16'h3e6a, 16'h494d,
// 16'h52b7, 16'h5a74, 16'h6057, 16'h644e,
// 16'h6635, 16'h660f, 16'h63d5, 16'h5f96,
// 16'h5966, 16'h5169, 16'h47c2, 16'h3ca9,
// 16'h3056, 16'h2303, 16'h1505, 16'h068c,
// 16'hf7fe, 16'he991, 16'hdb9d, 16'hce63,
// 16'hc22b, 16'hb735, 16'hadb8, 16'ha5e5,
// 16'h9fe8, 16'h9bd8, 16'h99d8, 16'h99e1,
// 16'h9c03, 16'ha027, 16'ha63f, 16'hae28,
// 16'hb7b8, 16'hc2c0, 16'hcf09, 16'hdc48,
// 16'hea4b, 16'hf8b5, 16'h0749, 16'h15ba,
// 16'h23b3, 16'h30fa, 16'h3d3f, 16'h4848,
// 16'h51d7, 16'h59c4, 16'h5fd5, 16'h6420,
// 16'h661d, 16'h6629, 16'h6428, 16'h6017,
// 16'h5a1d, 16'h5245, 16'h48cf, 16'h3dd1,
// 16'h319f, 16'h2463, 16'h166f, 16'h0802,
// 16'hf975, 16'heaf8, 16'hdd01, 16'hcfa6,
// 16'hc359, 16'hb83f, 16'hae95, 16'ha69c,
// 16'ha068, 16'h9c2b, 16'h99f3, 16'h99c9,
// 16'h9bb4, 16'h9fa6, 16'ha58e, 16'had49,
// 16'hb6b3, 16'hc196, 16'hcdc1, 16'hdaec,
// 16'he8de, 16'hf741, 16'h05d5, 16'h144b,
// 16'h2254, 16'h2fb2, 16'h3c11, 16'h473e,
// 16'h50f5, 16'h590c, 16'h5f50, 16'h63ad,
// 16'h65fe, 16'h6641, 16'h6472, 16'h6095,
// 16'h5acd, 16'h5321, 16'h49d3, 16'h3efa,
// 16'h32e4, 16'h25bf, 16'h17db, 16'h0976,
// 16'hfae8, 16'hec6b, 16'hde5b, 16'hd0f6,
// 16'hc483, 16'hb94d, 16'haf7b, 16'ha752,
// 16'ha0f3, 16'h9c80, 16'h9a13, 16'h99b6,
// 16'h9b6b, 16'h9f2b, 16'ha4e1, 16'hac6e,
// 16'hb5b0, 16'hc070, 16'hcc7d, 16'hd992,
// 16'he770, 16'hf5cf, 16'h045f, 16'h12dd,
// 16'h20f4, 16'h2e65, 16'h3ae2, 16'h462e,
// 16'h5012, 16'h584c, 16'h5ecc, 16'h634e,
// 16'h65df, 16'h664f, 16'h64b9, 16'h6110,
// 16'h5b75, 16'h53fb, 16'h4ad3, 16'h401f,
// 16'h3427, 16'h2719, 16'h1945, 16'h0aec,
// 16'hfc5b, 16'hedda, 16'hdfbe, 16'hd240,
// 16'hc5ba, 16'hba57, 16'hb068, 16'ha80c,
// 16'ha182, 16'h9cda, 16'h9a3a, 16'h99a7,
// 16'h9b28, 16'h9eb3, 16'ha439, 16'hab99,
// 16'hb4b1, 16'hbf4d, 16'hcb3a, 16'hd83a,
// 16'he606, 16'hf45c, 16'h02ea, 16'h116c,
// 16'h1f93, 16'h2d16, 16'h39af, 16'h451e,
// 16'h4f22, 16'h5793, 16'h5e37, 16'h62f4,
// 16'h65b5, 16'h6659, 16'h64fd, 16'h6181,
// 16'h5c1e, 16'h54cc, 16'h4bd2, 16'h413e,
// 16'h356a, 16'h286e, 16'h1ab1, 16'h0c5e,
// 16'hfdce, 16'hef4f, 16'he11d, 16'hd393,
// 16'hc6ec, 16'hbb6c, 16'hb153, 16'ha8d2,
// 16'ha210, 16'h9d3e, 16'h9a63, 16'h999e,
// 16'h9aeb, 16'h9e41, 16'ha396, 16'haac7,
// 16'hb3b5, 16'hbe2f, 16'hc9fb, 16'hd6e4,
// 16'he49b, 16'hf2ea, 16'h0174, 16'h0ffd,
// 16'h1e2f, 16'h2bc4, 16'h387a, 16'h4408,
// 16'h4e33, 16'h56d0, 16'h5da1, 16'h6293,
// 16'h6585, 16'h6661, 16'h6536, 16'h61f5,
// 16'h5cb9, 16'h55a2, 16'h4cc3, 16'h4264,
// 16'h36a0, 16'h29cb, 16'h1c13, 16'h0dd3,
// 16'hff45, 16'hf0bc, 16'he286, 16'hd4e1,
// 16'hc825, 16'hbc84, 16'hb243, 16'ha997,
// 16'ha2aa, 16'h9da0, 16'h9a97, 16'h9998,
// 16'h9ab2, 16'h9dd5, 16'ha2f7, 16'ha9fb,
// 16'hb2bd, 16'hbd12, 16'hc8c0, 16'hd58d,
// 16'he338, 16'hf174, 16'h2001, 16'h0e8a,
// 16'h1cc9, 16'h2a73, 16'h3740, 16'h42ee,
// 16'h4d44, 16'h5603, 16'h5d0a, 16'h622b,
// 16'h654f, 16'h6667, 16'h6569, 16'h6260,
// 16'h5d57, 16'h5668, 16'h4dbe, 16'h437a,
// 16'h37de, 16'h2b1c, 16'h1d7c, 16'h0f43,
// 16'h20bb, 16'hf22f, 16'he3e9, 16'hd639,
// 16'hc95c, 16'hbda1, 16'hb338, 16'haa61,
// 16'ha345, 16'h9e0b, 16'h9acd, 16'h999b,
// 16'h9a7c, 16'h9d6f, 16'ha25b, 16'ha935,
// 16'hb1c9, 16'hbbfa, 16'hc786, 16'hd43b,
// 16'he1d1, 16'hf005, 16'hfe89, 16'h0d1b,
// 16'h1b5f, 16'h2920, 16'h3603, 16'h41d2,
// 16'h4c4c, 16'h5537, 16'h5c6b, 16'h61be,
// 16'h6517, 16'h6661, 16'h659c, 16'h62c4,
// 16'h5dee, 16'h5730, 16'h4ead, 16'h4493,
// 16'h3913, 16'h2c70, 16'h1edf, 16'h10b7,
// 16'h022c, 16'hf3a6, 16'he54d, 16'hd792,
// 16'hca97, 16'hbec0, 16'hb431, 16'hab30,
// 16'ha3e7, 16'h9e79, 16'h9b09, 16'h99a2,
// 16'h9a4d, 16'h9d0d, 16'ha1c6, 16'ha871,
// 16'hb0da, 16'hbae4, 16'hc651, 16'hd2e9,
// 16'he06f, 16'hee91, 16'hfd18, 16'h0ba3,
// 16'h19fb, 16'h27c5, 16'h34c8, 16'h40b0,
// 16'h4b52, 16'h5464, 16'h5bca, 16'h614a,
// 16'h64da, 16'h6658, 16'h65c6, 16'h6327,
// 16'h5e7d, 16'h57f4, 16'h4f97, 16'h45ab,
// 16'h3a44, 16'h2dc2, 16'h2041, 16'h1225,
// 16'h03a7, 16'hf511, 16'he6bf, 16'hd8e3,
// 16'hcbdc, 16'hbfdf, 16'hb52e, 16'hac05,
// 16'ha48b, 16'h9eef, 16'h9b49, 16'h99ad,
// 16'h9a27, 16'h9cab, 16'ha13b, 16'ha7ae,
// 16'haff1, 16'hb9d2, 16'hc51d, 16'hd19c,
// 16'hdf0c, 16'hed22, 16'hfba2, 16'h0a30,
// 16'h1891, 16'h266d, 16'h3384, 16'h3f8f,
// 16'h4a51, 16'h5390, 16'h5b21, 16'h60d4,
// 16'h6496, 16'h6648, 16'h65f1, 16'h637a,
// 16'h5f14, 16'h58a8, 16'h5089, 16'h46b1,
// 16'h3b7f, 16'h2f07, 16'h21a8, 16'h1393,
// 16'h0519, 16'hf68a, 16'he824, 16'hda41,
// 16'hcd1e, 16'hc103, 16'hb631, 16'hacda,
// 16'ha538, 16'h9f67, 16'h9b90, 16'h99be,
// 16'h9a02, 16'h9c56, 16'ha0ac, 16'ha6f7,
// 16'haf07, 16'hb8c6, 16'hc3ec, 16'hd050,
// 16'hddab, 16'hebb5, 16'hfa2c, 16'h08bd,
// 16'h1724, 16'h2513, 16'h323f, 16'h3e6b,
// 16'h494c, 16'h52b8, 16'h5a71, 16'h605c,
// 16'h6448, 16'h663b, 16'h660b, 16'h63d6,
// 16'h5f98, 16'h5963, 16'h516b, 16'h47c0,
// 16'h3cac, 16'h3052, 16'h2308, 16'h1520,
// 16'h068f, 16'hf7ff, 16'he98d, 16'hdba1,
// 16'hce5f, 16'hc22f, 16'hb733, 16'hadb9,
// 16'ha5e4, 16'h9fe8, 16'h9bd9, 16'h99d7,
// 16'h99e2, 16'h9c03, 16'ha026, 16'ha640,
// 16'hae28, 16'hb7b7, 16'hc2c2, 16'hcf06,
// 16'hdc4c, 16'hea48, 16'hf8b5, 16'h074b,
// 16'h15b7, 16'h23b6, 16'h30f8, 16'h3d40,
// 16'h4847, 16'h51da, 16'h59bf, 16'h5fd9,
// 16'h63fe, 16'h661d, 16'h662c, 16'h6424,
// 16'h6019, 16'h5a1c, 16'h5246, 16'h48ce,
// 16'h3dd3, 16'h319c, 16'h2466, 16'h166c,
// 16'h0805, 16'hf971, 16'heafd, 16'hdcfd,
// 16'hcfa9, 16'hc357, 16'hb83f, 16'hae96,
// 16'ha69b, 16'ha06a, 16'h9c29, 16'h99f5,
// 16'h99c6, 16'h9bb6, 16'h9fa6, 16'ha58d,
// 16'had4b, 16'hb6af, 16'hc19a, 16'hcdbd,
// 16'hdaf1, 16'he8d9, 16'hf744, 16'h05d4,
// 16'h144b, 16'h2255, 16'h2fb1, 16'h3c11,
// 16'h473e, 16'h50f6, 16'h590b, 16'h5f52,
// 16'h63ab, 16'h65fe, 16'h6642, 16'h6470,
// 16'h6099, 16'h5ac9, 16'h5324, 16'h49d1,
// 16'h3efc, 16'h32e2, 16'h25c1, 16'h17d8,
// 16'h097b, 16'hfae3, 16'hec6f, 16'hde58,
// 16'hd0f7, 16'hc485, 16'hb94a, 16'haf7d,
// 16'ha751, 16'ha0f3, 16'h9c81, 16'h9a11,
// 16'h99b8, 16'h9b69, 16'h9f2d, 16'ha4df,
// 16'hac70, 16'hb5ad, 16'hc073, 16'hcc7a,
// 16'hd995, 16'he76f, 16'hf5ce, 16'h045f,
// 16'h12dd, 16'h20f5, 16'h2e65, 16'h3ae1,
// 16'h4630, 16'h500e, 16'h5851, 16'h5ec7,
// 16'h6354, 16'h65d9, 16'h6654, 16'h64b5,
// 16'h6113, 16'h5b73, 16'h53fd, 16'h4ad0,
// 16'h4022, 16'h3425, 16'h271a, 16'h1945,
// 16'h0aec, 16'hfc59, 16'heddf, 16'hdfb8,
// 16'hd246, 16'hc5b5, 16'hba5a, 16'hb066,
// 16'ha80e, 16'ha181, 16'h9cdb, 16'h9a39,
// 16'h99a7, 16'h9b28, 16'h9eb3, 16'ha43b,
// 16'hab96, 16'hb4b4, 16'hbf4a, 16'hcb3d,
// 16'hd837, 16'he609, 16'hf458, 16'h02ee,
// 16'h1169, 16'h1f95, 16'h2d15, 16'h39af,
// 16'h451d, 16'h4f25, 16'h5790, 16'h5e38,
// 16'h62f6, 16'h65b0, 16'h6660, 16'h64f7,
// 16'h6185, 16'h5c1b, 16'h54d0, 16'h4bcd,
// 16'h4144, 16'h3564, 16'h2872, 16'h1ab0,
// 16'h0c5d, 16'hfdd1, 16'hef4b, 16'he120,
// 16'hd391, 16'hc6ed, 16'hbb6c, 16'hb153,
// 16'ha8d0, 16'ha213, 16'h9d3b, 16'h9a66,
// 16'h999c, 16'h9aeb, 16'h9e41, 16'ha397,
// 16'haac5, 16'hb3b9, 16'hbe29, 16'hca01,
// 16'hd6de, 16'he4a0, 16'hf2e8, 16'h0174,
// 16'h0ffe, 16'h1e2c, 16'h2bc8, 16'h3877,
// 16'h4409, 16'h4e34, 16'h56ce, 16'h5da3,
// 16'h6292, 16'h6583, 16'h6665, 16'h6534,
// 16'h61f5, 16'h5cba, 16'h55a0, 16'h4cc5,
// 16'h4265, 16'h369d, 16'h29ce, 16'h1c11,
// 16'h0dd5, 16'hff43, 16'hf0be, 16'he283,
// 16'hd4e5, 16'hc821, 16'hbc87, 16'hb242,
// 16'ha997, 16'ha2aa, 16'h9d9f, 16'h9a98,
// 16'h9999, 16'h9ab0, 16'h9dd6, 16'ha2f6,
// 16'ha9fc, 16'hb2be, 16'hbd10, 16'hc8c2,
// 16'hd58b, 16'he339, 16'hf174, 16'h2001,
// 16'h0e8b, 16'h1cc7, 16'h2a75, 16'h373e,
// 16'h42f0, 16'h4d41, 16'h5606, 16'h5d08,
// 16'h622c, 16'h654e, 16'h6667, 16'h656a,
// 16'h625f, 16'h5d57, 16'h5669, 16'h4dbd,
// 16'h437a, 16'h37df, 16'h2b19, 16'h1d80,
// 16'h0f40, 16'h20bc, 16'hf230, 16'he3e7,
// 16'hd63a, 16'hc95c, 16'hbda0, 16'hb339,
// 16'haa62, 16'ha343, 16'h9e0c, 16'h9acd,
// 16'h999b, 16'h9a7d, 16'h9d6d, 16'ha25d,
// 16'ha934, 16'hb1c9, 16'hbbfb, 16'hc784,
// 16'hd43d, 16'he1d0, 16'hf005, 16'hfe8a,
// 16'h0d19, 16'h1b61, 16'h291e, 16'h3604,
// 16'h41d3, 16'h4c4a, 16'h5539, 16'h5c6a,
// 16'h61be, 16'h6517, 16'h6661, 16'h659d,
// 16'h62c2, 16'h5df1, 16'h572d, 16'h4eae,
// 16'h4494, 16'h3912, 16'h2c70, 16'h1ee0,
// 16'h10b4, 16'h0231, 16'hf3a0, 16'he553,
// 16'hd78d, 16'hca9b, 16'hbebd, 16'hb433,
// 16'hab2f, 16'ha3e7, 16'h9e7a, 16'h9b08,
// 16'h99a2, 16'h9a4f, 16'h9d09, 16'ha1cb,
// 16'ha86c, 16'hb0de, 16'hbae2, 16'hc651,
// 16'hd2eb, 16'he06a, 16'hee98, 16'hfd12,
// 16'h0ba7, 16'h19fa, 16'h27c4, 16'h34c8,
// 16'h40b1, 16'h4b50, 16'h5467, 16'h5bc8,
// 16'h614b, 16'h64d9, 16'h6658, 16'h65c7,
// 16'h6326, 16'h5e7e, 16'h57f4, 16'h4f97,
// 16'h45aa, 16'h3a45, 16'h2dc1, 16'h2042,
// 16'h1226, 16'h03a4, 16'hf515, 16'he6ba,
// 16'hd8e8, 16'hcbd9, 16'hbfe0, 16'hb52f,
// 16'hac03, 16'ha48c, 16'h9eef, 16'h9b48,
// 16'h99b0, 16'h9a23, 16'h9cae, 16'ha139,
// 16'ha7af, 16'haff2, 16'hb9cf, 16'hc520,
// 16'hd19a, 16'hdf0e, 16'hed20, 16'hfba4,
// 16'h0a2e, 16'h1893, 16'h266b, 16'h3386,
// 16'h3f8d, 16'h4a53, 16'h538f, 16'h5b21,
// 16'h60d4, 16'h6495, 16'h664a, 16'h65ee,
// 16'h637e, 16'h5f0f, 16'h58ad, 16'h5084,
// 16'h46b6, 16'h3b7a, 16'h2f0b, 16'h21a6,
// 16'h1393, 16'h051a, 16'hf68a, 16'he822,
// 16'hda44, 16'hcd1b, 16'hc105, 16'hb62f,
// 16'hacdd, 16'ha533, 16'h9f6d, 16'h9b8a,
// 16'h99c4, 16'h99fc, 16'h9c5a, 16'ha0ab,
// 16'ha6f6, 16'haf09, 16'hb8c4, 16'hc3ed,
// 16'hd052, 16'hdda8, 16'hebb6, 16'hfa2c,
// 16'h08bd, 16'h1725, 16'h2512, 16'h3240,
// 16'h3e68, 16'h494f, 16'h52b7, 16'h5a71,
// 16'h605c, 16'h644a, 16'h6636, 16'h6611,
// 16'h63d2, 16'h5f98, 16'h5966, 16'h5169,
// 16'h47c0, 16'h3cad, 16'h3050, 16'h230a,
// 16'h14ff, 16'h068f, 16'hf7ff, 16'he98e,
// 16'hdb9f, 16'hce62, 16'hc22b, 16'hb737,
// 16'hadb6, 16'ha5e5, 16'h9fe9, 16'h9bd7,
// 16'h99d9, 16'h99e1, 16'h9c01, 16'ha02a,
// 16'ha63d, 16'hae29, 16'hb7b8, 16'hc2c0,
// 16'hcf08, 16'hdc4a, 16'hea49, 16'hf8b6,
// 16'h0749, 16'h15b9, 16'h23b4, 16'h30fa,
// 16'h3d3e, 16'h4849, 16'h51d6, 16'h59c4,
// 16'h5fd7, 16'h63fe, 16'h661e, 16'h6628,
// 16'h6429, 16'h6017, 16'h5a1c, 16'h5247,
// 16'h48cc, 16'h3dd4, 16'h319e, 16'h2462,
// 16'h1670, 16'h0802, 16'hf973, 16'heafc,
// 16'hdcfd, 16'hcfa9, 16'hc358, 16'hb83d,
// 16'hae98, 16'ha69a, 16'ha06a, 16'h9c2a,
// 16'h99f2, 16'h99ca, 16'h9bb3, 16'h9fa9,
// 16'ha58a, 16'had4d, 16'hb6af, 16'hc198,
// 16'hcdc1, 16'hdaec, 16'he8df, 16'hf73e,
// 16'h05d9, 16'h1446, 16'h225a, 16'h2fad,
// 16'h3c14, 16'h473c, 16'h50f7, 16'h5909,
// 16'h5f55, 16'h63a8, 16'h6601, 16'h6640,
// 16'h6471, 16'h6099, 16'h5ac8, 16'h5325,
// 16'h49d0, 16'h3efd, 16'h32e2, 16'h25c0,
// 16'h17da, 16'h0978, 16'hfae6, 16'hec6b,
// 16'hde5c, 16'hd0f6, 16'hc484, 16'hb94c,
// 16'haf79, 16'ha755, 16'ha0f1, 16'h9c82,
// 16'h9a11, 16'h99b7, 16'h9b6a, 16'h9f2c,
// 16'ha4df, 16'hac70, 16'hb5b0, 16'hc06f,
// 16'hcc7d, 16'hd992, 16'he770, 16'hf5d0,
// 16'h045e, 16'h12de, 16'h20f3, 16'h2e67,
// 16'h3ade, 16'h4634, 16'h500a, 16'h5856,
// 16'h5ec3, 16'h6354, 16'h65db, 16'h6651,
// 16'h64b9, 16'h6111, 16'h5b72, 16'h53ff,
// 16'h4ace, 16'h4025, 16'h3421, 16'h271f,
// 16'h1940, 16'h0aee, 16'hfc5b, 16'hedda,
// 16'hdfbe, 16'hd241, 16'hc5b7, 16'hba5b,
// 16'hb064, 16'ha811, 16'ha17e, 16'h9cdc,
// 16'h9a3a, 16'h99a6, 16'h9b29, 16'h9eb3,
// 16'ha439, 16'hab9a, 16'hb4af, 16'hbf4e,
// 16'hcb3b, 16'hd839, 16'he607, 16'hf45b,
// 16'h02e9, 16'h116f, 16'h1f90, 16'h2d19,
// 16'h39ac, 16'h451f, 16'h4f23, 16'h5792,
// 16'h5e37, 16'h62f5, 16'h65b2, 16'h665d,
// 16'h64fa, 16'h6183, 16'h5c1d, 16'h54cd,
// 16'h4bd0, 16'h4141, 16'h3567, 16'h2871,
// 16'h1aae, 16'h0c60, 16'hfdce, 16'hef4f,
// 16'he11c, 16'hd394, 16'hc6ea, 16'hbb6f,
// 16'hb151, 16'ha8d2, 16'ha211, 16'h9d3c,
// 16'h9a65, 16'h999e, 16'h9ae8, 16'h9e44,
// 16'ha393, 16'haaca, 16'hb3b5, 16'hbe2c,
// 16'hc9fd, 16'hd6e1, 16'he4a0, 16'hf2e6,
// 16'h0176, 16'h0ffc, 16'h1e2e, 16'h2bc7,
// 16'h3877, 16'h4408, 16'h4e37, 16'h56ca,
// 16'h5da7, 16'h628e, 16'h6587, 16'h6662,
// 16'h6535, 16'h61f4, 16'h5cbc, 16'h559d,
// 16'h4cc9, 16'h4260, 16'h36a2, 16'h29ca,
// 16'h1c13, 16'h0dd4, 16'hff43, 16'hf0c0,
// 16'he280, 16'hd4e7, 16'hc820, 16'hbc86,
// 16'hb244, 16'ha995, 16'ha2ac, 16'h9d9e,
// 16'h9a98, 16'h9998, 16'h9ab3, 16'h9dd3,
// 16'ha2f8, 16'ha9fb, 16'hb2be, 16'hbd11,
// 16'hc8c1, 16'hd58b, 16'he33a, 16'hf173,
// 16'h2002, 16'h0e89, 16'h1cc9, 16'h2a74,
// 16'h373f, 16'h42ef, 16'h4d42, 16'h5604,
// 16'h5d0a, 16'h622b, 16'h654f, 16'h6667,
// 16'h6569, 16'h625f, 16'h5d58, 16'h5669,
// 16'h4dbc, 16'h437c, 16'h37dc, 16'h2b1d,
// 16'h1d7c, 16'h0f43, 16'h20ba, 16'hf230,
// 16'he3e9, 16'hd638, 16'hc95e, 16'hbd9e,
// 16'hb33a, 16'haa61, 16'ha345, 16'h9e0c,
// 16'h9acb, 16'h999d, 16'h9a7b, 16'h9d6f,
// 16'ha25c, 16'ha934, 16'hb1ca, 16'hbbfa,
// 16'hc783, 16'hd440, 16'he1cc, 16'hf009,
// 16'hfe87, 16'h0d1a, 16'h1b62, 16'h291d,
// 16'h3606, 16'h41d0, 16'h4c4d, 16'h5536,
// 16'h5c6c, 16'h61be, 16'h6517, 16'h6661,
// 16'h659c, 16'h62c4, 16'h5ded, 16'h5731,
// 16'h4eac, 16'h4494, 16'h3914, 16'h2c6e,
// 16'h1ee1, 16'h10b4, 16'h022f, 16'hf3a4,
// 16'he54f, 16'hd791, 16'hca98, 16'hbebe,
// 16'hb432, 16'hab31, 16'ha3e6, 16'h9e7a,
// 16'h9b09, 16'h999f, 16'h9a52, 16'h9d08,
// 16'ha1cb, 16'ha86c, 16'hb0de, 16'hbae2,
// 16'hc651, 16'hd2ea, 16'he06d, 16'hee94,
// 16'hfd15, 16'h0ba6, 16'h19f7, 16'h27cb,
// 16'h34c1, 16'h40b5, 16'h4b50, 16'h5464,
// 16'h5bcb, 16'h6149, 16'h64da, 16'h6659,
// 16'h65c5, 16'h6327, 16'h5e7d, 16'h57f4,
// 16'h4f99, 16'h45a7, 16'h3a48, 16'h2dbe,
// 16'h2044, 16'h1224, 16'h03a6, 16'hf514,
// 16'he6bb, 16'hd8e6, 16'hcbdb, 16'hbfde,
// 16'hb531, 16'hac01, 16'ha48e, 16'h9eee,
// 16'h9b48, 16'h99b0, 16'h9a23, 16'h9caf,
// 16'ha138, 16'ha7af, 16'haff2, 16'hb9d0,
// 16'hc51f, 16'hd19b, 16'hdf0b, 16'hed24,
// 16'hfb9f, 16'h0a34, 16'h188e, 16'h266e,
// 16'h3384, 16'h3f8f, 16'h4a50, 16'h5393,
// 16'h5b1d, 16'h60d8, 16'h6493, 16'h664a,
// 16'h65ee, 16'h637f, 16'h5f0e, 16'h58ae,
// 16'h5083, 16'h46b6, 16'h3b7c, 16'h2f09,
// 16'h21a6, 16'h1394, 16'h0519, 16'hf689,
// 16'he826, 16'hda3f, 16'hcd1f, 16'hc102,
// 16'hb632, 16'hacd9, 16'ha539, 16'h9f66,
// 16'h9b90, 16'h99c0, 16'h9a20, 16'h9c56,
// 16'ha0ad, 16'ha6f5, 16'haf0b, 16'hb8c2,
// 16'hc3ef, 16'hd04f, 16'hddaa, 16'hebb6,
// 16'hfa2b, 16'h08bd, 16'h1726, 16'h2511,
// 16'h3241, 16'h3e68, 16'h494e, 16'h52b6,
// 16'h5a74, 16'h6059, 16'h644c, 16'h6636,
// 16'h660f, 16'h63d4, 16'h5f97, 16'h5967,
// 16'h5167, 16'h47c3, 16'h3caa, 16'h3052,
// 16'h230a, 16'h14fd, 16'h0693, 16'hf7fa,
// 16'he993, 16'hdb9a, 16'hce65, 16'hc22c,
// 16'hb733, 16'hadba, 16'ha5e3, 16'h9fe7,
// 16'h9bdd, 16'h99d2, 16'h99e7, 16'h9bfd,
// 16'ha02c, 16'ha63b, 16'hae2c, 16'hb7b4,
// 16'hc2c5, 16'hcf03, 16'hdc4e, 16'hea47,
// 16'hf8b5, 16'h074c, 16'h15b6, 16'h23b7,
// 16'h30f8, 16'h3d3e, 16'h4849, 16'h51d8,
// 16'h59c1, 16'h5fd9, 16'h63fd, 16'h661e,
// 16'h662a, 16'h6426, 16'h6019, 16'h5a1b,
// 16'h5247, 16'h48cd, 16'h3dd3, 16'h319e,
// 16'h2463, 16'h166e, 16'h0804, 16'hf971,
// 16'heafe, 16'hdcfc, 16'hcfa9, 16'hc358,
// 16'hb83d, 16'hae99, 16'ha699, 16'ha069,
// 16'h9c2c, 16'h99f0, 16'h99cc, 16'h9bb3,
// 16'h9fa5, 16'ha590, 16'had47, 16'hb6b3,
// 16'hc197, 16'hcdc0, 16'hdaed, 16'he8de,
// 16'hf73f, 16'h05d7, 16'h144a, 16'h2256,
// 16'h2faf, 16'h3c13, 16'h473d, 16'h50f5,
// 16'h590e, 16'h5f4e, 16'h63af, 16'h65fc,
// 16'h6643, 16'h646f, 16'h609a, 16'h5ac7,
// 16'h5327, 16'h49cf, 16'h3efc, 16'h32e3,
// 16'h25bf, 16'h17db, 16'h0978, 16'hfae5,
// 16'hec6e, 16'hde58, 16'hd0f8, 16'hc483,
// 16'hb94c, 16'haf7c, 16'ha751, 16'ha0f3,
// 16'h9c81, 16'h9a11, 16'h99b9, 16'h9b67,
// 16'h9f2e, 16'ha4de, 16'hac71, 16'hb5af,
// 16'hc070, 16'hcc7c, 16'hd993, 16'he770,
// 16'hf5ce, 16'h0461, 16'h12da, 16'h20f7,
// 16'h2e64, 16'h3ae1, 16'h4630, 16'h500e,
// 16'h5852, 16'h5ec6, 16'h6354, 16'h65d9,
// 16'h6654, 16'h64b6, 16'h6112, 16'h5b73,
// 16'h53fd, 16'h4ad1, 16'h4021, 16'h3425,
// 16'h271a, 16'h1945, 16'h0aec, 16'hfc5a,
// 16'heddd, 16'hdfba, 16'hd245, 16'hc5b5,
// 16'hba5a, 16'hb067, 16'ha80c, 16'ha184,
// 16'h9cd8, 16'h9a3b, 16'h99a7, 16'h9b25,
// 16'h9eb9, 16'ha433, 16'hab9e, 16'hb4ae,
// 16'hbf4d, 16'hcb3c, 16'hd838, 16'he607,
// 16'hf45b, 16'h02ea, 16'h116e, 16'h1f90,
// 16'h2d19, 16'h39ac, 16'h4520, 16'h4f22,
// 16'h5792, 16'h5e38, 16'h62f4, 16'h65b3,
// 16'h665c, 16'h64fa, 16'h6184, 16'h5c1c,
// 16'h54cd, 16'h4bd0, 16'h4142, 16'h3565,
// 16'h2874, 16'h1aab, 16'h0c62, 16'hfdcd,
// 16'hef4f, 16'he11c, 16'hd394, 16'hc6eb,
// 16'hbb6d, 16'hb153, 16'ha8d0, 16'ha212,
// 16'h9d3c, 16'h9a65, 16'h999d, 16'h9aeb,
// 16'h9e40, 16'ha398, 16'haac5, 16'hb3b7,
// 16'hbe2d, 16'hc9fc, 16'hd6e3, 16'he49d,
// 16'hf2e9, 16'h0173, 16'h0fff, 16'h1e2c,
// 16'h2bc7, 16'h3879, 16'h4406, 16'h4e38,
// 16'h56ca, 16'h5da6, 16'h6290, 16'h6584,
// 16'h6666, 16'h6531, 16'h61f9, 16'h5cb6,
// 16'h55a3, 16'h4cc3, 16'h4265, 16'h369f,
// 16'h29cc, 16'h1c12, 16'h0dd4, 16'hff43,
// 16'hf0c0, 16'he281, 16'hd4e6, 16'hc820,
// 16'hbc88, 16'hb241, 16'ha999, 16'ha2a7,
// 16'h9da2, 16'h9a96, 16'h999a, 16'h9ab0,
// 16'h9dd6, 16'ha2f6, 16'ha9fc, 16'hb2bd,
// 16'hbd12, 16'hc8c0, 16'hd58d, 16'he338,
// 16'hf173, 16'h2003, 16'h0e88, 16'h1ccb,
// 16'h2a72, 16'h373f, 16'h42f0, 16'h4d41,
// 16'h5606, 16'h5d08, 16'h622c, 16'h654d,
// 16'h6669, 16'h6568, 16'h6261, 16'h5d55,
// 16'h566b, 16'h4db9, 16'h4381, 16'h37d7,
// 16'h2b22, 16'h1d77, 16'h0f46, 16'h20ba,
// 16'hf22e, 16'he3ec, 16'hd635, 16'hc960,
// 16'hbd9e, 16'hb339, 16'haa61, 16'ha346,
// 16'h9e0a, 16'h9ace, 16'h999a, 16'h9a7d,
// 16'h9d6e, 16'ha25c, 16'ha934, 16'hb1ca,
// 16'hbbf9, 16'hc787, 16'hd439, 16'he1d4,
// 16'hf001, 16'hfe8e, 16'h0d16, 16'h1b62,
// 16'h291f, 16'h3602, 16'h41d5, 16'h4c49,
// 16'h5539, 16'h5c6a, 16'h61be, 16'h6517,
// 16'h6662, 16'h659b, 16'h62c5, 16'h5ded,
// 16'h5731, 16'h4eab, 16'h4496, 16'h3911,
// 16'h2c70, 16'h1ee1, 16'h10b2, 16'h0234,
// 16'hf39d, 16'he555, 16'hd78c, 16'hca9c,
// 16'hbebd, 16'hb431, 16'hab32, 16'ha3e5,
// 16'h9e7b, 16'h9b08, 16'h99a1, 16'h9a4f,
// 16'h9d0c, 16'ha1c6, 16'ha871, 16'hb0da,
// 16'hbae5, 16'hc64f, 16'hd2ec, 16'he06a,
// 16'hee98, 16'hfd11, 16'h0ba8, 16'h19f9,
// 16'h27c6, 16'h34c6, 16'h40b2, 16'h4b50,
// 16'h5467, 16'h5bc7, 16'h614d, 16'h64d7,
// 16'h665a, 16'h65c6, 16'h6325, 16'h5e7f,
// 16'h57f3, 16'h4f98, 16'h45a9, 16'h3a47,
// 16'h2dbe, 16'h2045, 16'h1221, 16'h03aa,
// 16'hf510, 16'he6bf, 16'hd8e3, 16'hcbdc,
// 16'hbfdf, 16'hb52e, 16'hac05, 16'ha48b,
// 16'h9eef, 16'h9b49, 16'h99ae, 16'h9a24,
// 16'h9cb0, 16'ha135, 16'ha7b3, 16'hafee,
// 16'hb9d4, 16'hc51b, 16'hd19f, 16'hdf07,
// 16'hed27, 16'hfb9f, 16'h0a32, 16'h1891,
// 16'h266a, 16'h3388, 16'h3f8c, 16'h4a54,
// 16'h538f, 16'h5b20, 16'h60d5, 16'h6495,
// 16'h664a, 16'h65ee, 16'h637e, 16'h5f0f,
// 16'h58ad, 16'h5084, 16'h46b6, 16'h3b7a,
// 16'h2f0b, 16'h21a6, 16'h1393, 16'h051b,
// 16'hf687, 16'he827, 16'hda3f, 16'hcd1f,
// 16'hc102, 16'hb631, 16'hacdb, 16'ha536,
// 16'h9f69, 16'h9b8e, 16'h99c0, 16'h9a20,
// 16'h9c56, 16'ha0ad, 16'ha6f6, 16'haf0a,
// 16'hb8c1, 16'hc3f1, 16'hd04d, 16'hddac,
// 16'hebb5, 16'hfa2b, 16'h08be, 16'h1725,
// 16'h2511, 16'h3240, 16'h3e6a, 16'h494d,
// 16'h52b7, 16'h5a74, 16'h6056, 16'h6450,
// 16'h6633, 16'h6611, 16'h63d3, 16'h5f97,
// 16'h5967, 16'h5167, 16'h47c3, 16'h3ca9,
// 16'h3055, 16'h2306, 16'h1501, 16'h068f,
// 16'hf7fc, 16'he993, 16'hdb9b, 16'hce64,
// 16'hc22b, 16'hb735, 16'hadb7, 16'ha5e7,
// 16'h9fe5, 16'h9bdc, 16'h99d4, 16'h99e4,
// 16'h9c01, 16'ha028, 16'ha640, 16'hae26,
// 16'hb7b9, 16'hc2c2, 16'hcf04, 16'hdc4f,
// 16'hea45, 16'hf8b8, 16'h0749, 16'h15b8,
// 16'h23b5, 16'h30fa, 16'h3d3e, 16'h4848,
// 16'h51d8, 16'h59c1, 16'h5fda, 16'h63fc,
// 16'h661f, 16'h6628, 16'h6427, 16'h601a,
// 16'h5a19, 16'h524a, 16'h48c9, 16'h3dd7,
// 16'h319a, 16'h2467, 16'h166b, 16'h0807,
// 16'hf96e, 16'heb02, 16'hdcf6, 16'hcfb0,
// 16'hc351, 16'hb844, 16'hae93, 16'ha69c,
// 16'ha069, 16'h9c2b, 16'h99f1, 16'h99cb,
// 16'h9bb2, 16'h9fa9, 16'ha58c, 16'had49,
// 16'hb6b2, 16'hc198, 16'hcdbf, 16'hdaf0,
// 16'he8d9, 16'hf743, 16'h05d6, 16'h1449,
// 16'h2257, 16'h2fb0, 16'h3c11, 16'h473f,
// 16'h50f4, 16'h590c, 16'h5f52, 16'h63ab,
// 16'h65ff, 16'h6641, 16'h6470, 16'h6099,
// 16'h5ac9, 16'h5324, 16'h49d2, 16'h3efa,
// 16'h32e4, 16'h25bf, 16'h17da, 16'h0979,
// 16'hfae5, 16'hec6d, 16'hde59, 16'hd0f7,
// 16'hc483, 16'hb94e, 16'haf79, 16'ha753,
// 16'ha0f3, 16'h9c7f, 16'h9a15, 16'h99b4,
// 16'h9b6c, 16'h9f2a, 16'ha4e2, 16'hac6e,
// 16'hb5b0, 16'hc06f, 16'hcc7e, 16'hd991,
// 16'he772, 16'hf5cd, 16'h0460, 16'h12dc,
// 16'h20f6, 16'h2e62, 16'h3ae6, 16'h462a,
// 16'h5013, 16'h584f, 16'h5ec6, 16'h6356,
// 16'h65d7, 16'h6655, 16'h64b5, 16'h6113,
// 16'h5b73, 16'h53fe, 16'h4ace, 16'h4025,
// 16'h3421, 16'h271e, 16'h1942, 16'h0aed,
// 16'hfc5b, 16'heddb, 16'hdfbc, 16'hd243,
// 16'hc5b6, 16'hba5c, 16'hb063, 16'ha811,
// 16'ha17e, 16'h9cdd, 16'h9a38, 16'h99a9,
// 16'h9b26, 16'h9eb5, 16'ha437, 16'hab9b,
// 16'hb4af, 16'hbf4f, 16'hcb39, 16'hd83a,
// 16'he607, 16'hf45a, 16'h02ec, 16'h116a,
// 16'h1f95, 16'h2d15, 16'h39af, 16'h451e,
// 16'h4f22, 16'h5793, 16'h5e37, 16'h62f5,
// 16'h65b1, 16'h6660, 16'h64f5, 16'h6189,
// 16'h5c18, 16'h54d0, 16'h4bcf, 16'h4141,
// 16'h3568, 16'h286f, 16'h1ab1, 16'h0c5d,
// 16'hfdcf, 16'hef50, 16'he11a, 16'hd396,
// 16'hc6e8, 16'hbb70, 16'hb151, 16'ha8d2,
// 16'ha211, 16'h9d3c, 16'h9a64, 16'h999f,
// 16'h9ae8, 16'h9e44, 16'ha394, 16'haac8,
// 16'hb3b6, 16'hbe2c, 16'hc9fd, 16'hd6e2,
// 16'he49e, 16'hf2e8, 16'h0176, 16'h0ffa,
// 16'h1e30, 16'h2bc5, 16'h3879, 16'h4408,
// 16'h4e36, 16'h56cc, 16'h5da3, 16'h6293,
// 16'h6583, 16'h6665, 16'h6534, 16'h61f4,
// 16'h5cbc, 16'h559d, 16'h4cca, 16'h425e,
// 16'h36a4, 16'h29c8, 16'h1c15, 16'h0dd2,
// 16'hff47, 16'hf0ba, 16'he285, 16'hd4e3,
// 16'hc823, 16'hbc86, 16'hb243, 16'ha996,
// 16'ha2a9, 16'h9da2, 16'h9a95, 16'h999b,
// 16'h9ab0, 16'h9dd5, 16'ha2f6, 16'ha9fe,
// 16'hb2ba, 16'hbd15, 16'hc8bd, 16'hd58f,
// 16'he337, 16'hf175, 16'h2020, 16'h0e8b,
// 16'h1cc8, 16'h2a74, 16'h373f, 16'h42f0,
// 16'h4d40, 16'h5607, 16'h5d08, 16'h622b,
// 16'h6550, 16'h6665, 16'h656a, 16'h6261,
// 16'h5d54, 16'h566d, 16'h4db8, 16'h4380,
// 16'h37d8, 16'h2b21, 16'h1d78, 16'h0f47,
// 16'h20b8, 16'hf230, 16'he3e9, 16'hd639,
// 16'hc95d, 16'hbd9f, 16'hb339, 16'haa61,
// 16'ha345, 16'h9e0d, 16'h9ac9, 16'h999f,
// 16'h9a79, 16'h9d70, 16'ha25c, 16'ha933,
// 16'hb1cc, 16'hbbf7, 16'hc788, 16'hd439,
// 16'he1d3, 16'hf003, 16'hfe8d, 16'h0d14,
// 16'h1b66, 16'h291b, 16'h3606, 16'h41d2,
// 16'h4c4a, 16'h5538, 16'h5c6c, 16'h61bc,
// 16'h6519, 16'h6660, 16'h659c, 16'h62c4,
// 16'h5dee, 16'h572f, 16'h4eaf, 16'h4491,
// 16'h3915, 16'h2c6e, 16'h1ee1, 16'h10b4,
// 16'h0230, 16'hf3a2, 16'he550, 16'hd791,
// 16'hca97, 16'hbec0, 16'hb431, 16'hab30,
// 16'ha3e7, 16'h9e79, 16'h9b0a, 16'h999f,
// 16'h9a51, 16'h9d0a, 16'ha1c7, 16'ha872,
// 16'hb0d8, 16'hbae6, 16'hc650, 16'hd2e9,
// 16'he06e, 16'hee94, 16'hfd15, 16'h0ba5,
// 16'h19fa, 16'h27c6, 16'h34c6, 16'h40b2,
// 16'h4b50, 16'h5467, 16'h5bc8, 16'h614a,
// 16'h64db, 16'h6655, 16'h65cc, 16'h6320,
// 16'h5e83, 16'h57ef, 16'h4f9d, 16'h45a3,
// 16'h3a4d, 16'h2db8, 16'h204a, 16'h121f,
// 16'h03aa, 16'hf511, 16'he6bd, 16'hd8e5,
// 16'hcbdb, 16'hbfdf, 16'hb52e, 16'hac07,
// 16'ha488, 16'h9ef2, 16'h9b46, 16'h99af,
// 16'h9a26, 16'h9cac, 16'ha13b, 16'ha7ad,
// 16'haff2, 16'hb9d1, 16'hc51d, 16'hd19e,
// 16'hdf09, 16'hed25, 16'hfba0, 16'h0a31,
// 16'h1890, 16'h266e, 16'h3383, 16'h3f91,
// 16'h4a4f, 16'h5392, 16'h5b1f, 16'h60d6,
// 16'h6493, 16'h664d, 16'h65ea, 16'h6383,
// 16'h5f0a, 16'h58b1, 16'h5081, 16'h46b8,
// 16'h3b79, 16'h2f0b, 16'h21a6, 16'h1393,
// 16'h051c, 16'hf685, 16'he829, 16'hda3d,
// 16'hcd20, 16'hc103, 16'hb62f, 16'hacdd,
// 16'ha536, 16'h9f67, 16'h9b91, 16'h99bc,
// 16'h9a04, 16'h9c55, 16'ha0ac, 16'ha6f7,
// 16'haf07, 16'hb8c7, 16'hc3ea, 16'hd054,
// 16'hdda6, 16'hebb9, 16'hfa28, 16'h08c1,
// 16'h1722, 16'h2515, 16'h323d, 16'h3e6b,
// 16'h494c, 16'h52b9, 16'h5a71, 16'h605b,
// 16'h644b, 16'h6636, 16'h6610, 16'h63d3,
// 16'h5f98, 16'h5966, 16'h5167, 16'h47c4,
// 16'h3ca8, 16'h3056, 16'h2304, 16'h1502,
// 16'h0690, 16'hf7fc, 16'he992, 16'hdb9a,
// 16'hce65, 16'hc22b, 16'hb736, 16'hadb6,
// 16'ha5e7, 16'h9fe5, 16'h9bdc, 16'h99d5,
// 16'h99e2, 16'h9c03, 16'ha027, 16'ha63f,
// 16'hae28, 16'hb7b8, 16'hc2c1, 16'hcf07,
// 16'hdc4a, 16'hea4a, 16'hf8b4, 16'h074c,
// 16'h15b6, 16'h23b6, 16'h30fa, 16'h3d3d,
// 16'h484a, 16'h51d5, 16'h59c5, 16'h5fd5,
// 16'h6401, 16'h661b, 16'h662c, 16'h6424,
// 16'h601b, 16'h5a19, 16'h5249, 16'h48cd,
// 16'h3dd1, 16'h31a1, 16'h2460, 16'h1670,
// 16'h0804, 16'hf970, 16'heaff, 16'hdcfb,
// 16'hcfaa, 16'hc357, 16'hb83f, 16'hae95,
// 16'ha69e, 16'ha064, 16'h9c31, 16'h99ec,
// 16'h99ce, 16'h9bb1, 16'h9fa9, 16'ha58b,
// 16'had4b, 16'hb6b0, 16'hc19a, 16'hcdbd,
// 16'hdaf1, 16'he8d9, 16'hf743, 16'h05d5,
// 16'h144b, 16'h2255, 16'h2fb1, 16'h3c11,
// 16'h473d, 16'h50f7, 16'h590a, 16'h5f53,
// 16'h63ab, 16'h65fe, 16'h6642, 16'h646f,
// 16'h609a, 16'h5ac8, 16'h5326, 16'h49cf,
// 16'h3efd, 16'h32e2, 16'h25bf, 16'h17dc,
// 16'h0977, 16'hfae6, 16'hec6c, 16'hde5b,
// 16'hd0f5, 16'hc486, 16'hb949, 16'haf7d,
// 16'ha752, 16'ha0f3, 16'h9c80, 16'h9a12,
// 16'h99b7, 16'h9b6a, 16'h9f2c, 16'ha4e0,
// 16'hac6f, 16'hb5af, 16'hc071, 16'hcc7c,
// 16'hd992, 16'he771, 16'hf5ce, 16'h045f,
// 16'h12de, 16'h20f3, 16'h2e66, 16'h3ae1,
// 16'h462f, 16'h5010, 16'h584f, 16'h5ec9,
// 16'h6352, 16'h65db, 16'h6652, 16'h64b7,
// 16'h6110, 16'h5b78, 16'h53f7, 16'h4ad6,
// 16'h401d, 16'h3428, 16'h2719, 16'h1944,
// 16'h0aee, 16'hfc58, 16'hedde, 16'hdfba,
// 16'hd243, 16'hc5b8, 16'hba59, 16'hb065,
// 16'ha80f, 16'ha180, 16'h9cdb, 16'h9a3a,
// 16'h99a7, 16'h9b27, 16'h9eb4, 16'ha439,
// 16'hab98, 16'hb4b3, 16'hbf4b, 16'hcb3c,
// 16'hd839, 16'he606, 16'hf45b, 16'h02ec,
// 16'h116a, 16'h1f96, 16'h2d12, 16'h39b2,
// 16'h451c, 16'h4f24, 16'h5792, 16'h5e36,
// 16'h62f7, 16'h65b0, 16'h665f, 16'h64f7,
// 16'h6187, 16'h5c19, 16'h54d0, 16'h4bce,
// 16'h4142, 16'h3566, 16'h2873, 16'h1aac,
// 16'h0c61, 16'hfdce, 16'hef4e, 16'he11d,
// 16'hd394, 16'hc6e9, 16'hbb70, 16'hb151,
// 16'ha8d1, 16'ha213, 16'h9d3a, 16'h9a66,
// 16'h999e, 16'h9ae8, 16'h9e44, 16'ha394,
// 16'haac8, 16'hb3b6, 16'hbe2d, 16'hc9fb,
// 16'hd6e4, 16'he49c, 16'hf2e9, 16'h0176,
// 16'h0ffa, 16'h1e31, 16'h2bc3, 16'h387b,
// 16'h4406, 16'h4e37, 16'h56cc, 16'h5da3,
// 16'h6293, 16'h6582, 16'h6666, 16'h6532,
// 16'h61f7, 16'h5cba, 16'h559e, 16'h4cc8,
// 16'h4260, 16'h36a3, 16'h29c9, 16'h1c15,
// 16'h0dd2, 16'hff45, 16'hf0bd, 16'he284,
// 16'hd4e3, 16'hc824, 16'hbc84, 16'hb244,
// 16'ha997, 16'ha2a8, 16'h9da2, 16'h9a95,
// 16'h999a, 16'h9ab2, 16'h9dd3, 16'ha2f9,
// 16'ha9f8, 16'hb2c1, 16'hbd0f, 16'hc8c2,
// 16'hd58c, 16'he337, 16'hf176, 16'h2020,
// 16'h0e89, 16'h1ccb, 16'h2a72, 16'h3740,
// 16'h42ee, 16'h4d43, 16'h5603, 16'h5d0c,
// 16'h6229, 16'h6550, 16'h6665, 16'h656c,
// 16'h625d, 16'h5d5a, 16'h5666, 16'h4dbe,
// 16'h437c, 16'h37db, 16'h2b1f, 16'h1d79,
// 16'h0f46, 16'h20b9, 16'hf22f, 16'he3ea,
// 16'hd638, 16'hc95d, 16'hbda0, 16'hb338,
// 16'haa62, 16'ha345, 16'h9e0a, 16'h9ace,
// 16'h999a, 16'h9a7e, 16'h9d6c, 16'ha25f,
// 16'ha930, 16'hb1ce, 16'hbbf6, 16'hc787,
// 16'hd43d, 16'he1cd, 16'hf008, 16'hfe88,
// 16'h0d1a, 16'h1b62, 16'h291c, 16'h3606,
// 16'h41d1, 16'h4c4d, 16'h5536, 16'h5c6c,
// 16'h61bd, 16'h6518, 16'h6660, 16'h659e,
// 16'h62c1, 16'h5df1, 16'h572d, 16'h4eb0,
// 16'h4490, 16'h3917, 16'h2c6b, 16'h1ee4,
// 16'h10b2, 16'h0231, 16'hf3a2, 16'he550,
// 16'hd790, 16'hca99, 16'hbebe, 16'hb432,
// 16'hab30, 16'ha3e7, 16'h9e79, 16'h9b09,
// 16'h99a1, 16'h9a50, 16'h9d09, 16'ha1ca,
// 16'ha86d, 16'hb0dd, 16'hbae4, 16'hc64f,
// 16'hd2ec, 16'he06b, 16'hee95, 16'hfd15,
// 16'h0ba6, 16'h19f8, 16'h27c9, 16'h34c2,
// 16'h40b5, 16'h4b4f, 16'h5466, 16'h5bca,
// 16'h6149, 16'h64db, 16'h6656, 16'h65c9,
// 16'h6324, 16'h5e80, 16'h57f1, 16'h4f9b,
// 16'h45a5, 16'h3a4b, 16'h2dbc, 16'h2044,
// 16'h1225, 16'h03a4, 16'hf516, 16'he6ba,
// 16'hd8e6, 16'hcbdc, 16'hbfdc, 16'hb532,
// 16'hac01, 16'ha48f, 16'h9eeb, 16'h9b4d,
// 16'h99a9, 16'h9a29, 16'h9cac, 16'ha139,
// 16'ha7af, 16'haff2, 16'hb9cf, 16'hc520,
// 16'hd19b, 16'hdf0b, 16'hed24, 16'hfba0,
// 16'h0a32, 16'h188f, 16'h266e, 16'h3385,
// 16'h3f8c, 16'h4a56, 16'h538b, 16'h5b25,
// 16'h60d1, 16'h6497, 16'h664a, 16'h65ed,
// 16'h6380, 16'h5f0d, 16'h58af, 16'h5082,
// 16'h46b8, 16'h3b79, 16'h2f0c, 16'h21a4,
// 16'h1394, 16'h051b, 16'hf687, 16'he827,
// 16'hda3e, 16'hcd1f, 16'hc103, 16'hb631,
// 16'hacda, 16'ha538, 16'h9f67, 16'h9b90,
// 16'h99bd, 16'h9a04, 16'h9c52, 16'ha0b2,
// 16'ha6f0, 16'haf0f, 16'hb8be, 16'hc3f2,
// 16'hd04d, 16'hddab, 16'hebb7, 16'hfa28,
// 16'h08c1, 16'h1722, 16'h2513, 16'h3240,
// 16'h3e69, 16'h494e, 16'h52b6, 16'h5a74,
// 16'h6057, 16'h644e, 16'h6636, 16'h660e,
// 16'h63d6, 16'h5f95, 16'h5967, 16'h5168,
// 16'h47c3, 16'h3ca8, 16'h3056, 16'h2305,
// 16'h1502, 16'h068e, 16'hf7fe, 16'he990,
// 16'hdb9d, 16'hce63, 16'hc22b, 16'hb735,
// 16'hadb9, 16'ha5e3, 16'h9fe9, 16'h9bd9,
// 16'h99d6, 16'h99e4, 16'h9c20, 16'ha029,
// 16'ha63e, 16'hae28, 16'hb7b9, 16'hc2c0,
// 16'hcf08, 16'hdc49, 16'hea4a, 16'hf8b4,
// 16'h074d, 16'h15b4, 16'h23b9, 16'h30f6,
// 16'h3d41, 16'h4846, 16'h51da, 16'h59c0,
// 16'h5fda, 16'h63fc, 16'h661e, 16'h662b,
// 16'h6425, 16'h601b, 16'h5a18, 16'h524a,
// 16'h48ca, 16'h3dd6, 16'h319c, 16'h2465,
// 16'h166c, 16'h0807, 16'hf96d, 16'heb02,
// 16'hdcf8, 16'hcfad, 16'hc356, 16'hb83d,
// 16'hae99, 16'ha699, 16'ha069, 16'h9c2d,
// 16'h99ee, 16'h99ce, 16'h9bb0, 16'h9fab,
// 16'ha588, 16'had4e, 16'hb6ae, 16'hc19b,
// 16'hcdbc, 16'hdaf1, 16'he8da, 16'hf743,
// 16'h05d4, 16'h144a, 16'h2257, 16'h2faf,
// 16'h3c14, 16'h473b, 16'h50f7, 16'h590b,
// 16'h5f52, 16'h63ab, 16'h65ff, 16'h6641,
// 16'h6471, 16'h6097, 16'h5acb, 16'h5323,
// 16'h49d2, 16'h3efa, 16'h32e5, 16'h25bd,
// 16'h17dd, 16'h0975, 16'hfae9, 16'hec69,
// 16'hde5e, 16'hd0f2, 16'hc487, 16'hb94a,
// 16'haf7c, 16'ha752, 16'ha0f2, 16'h9c81,
// 16'h9a13, 16'h99b5, 16'h9b6b, 16'h9f2b,
// 16'ha4e1, 16'hac6e, 16'hb5b1, 16'hc06e,
// 16'hcc7e, 16'hd993, 16'he76e, 16'hf5d1,
// 16'h045e, 16'h12dd, 16'h20f5, 16'h2e64,
// 16'h3ae2, 16'h4630, 16'h500e, 16'h5851,
// 16'h5ec7, 16'h6353, 16'h65db, 16'h6651,
// 16'h64b8, 16'h6111, 16'h5b74, 16'h53fc,
// 16'h4ad2, 16'h401f, 16'h3428, 16'h2717,
// 16'h1948, 16'h0ae9, 16'hfc5c, 16'heddc,
// 16'hdfba, 16'hd245, 16'hc5b6, 16'hba59,
// 16'hb067, 16'ha80d, 16'ha182, 16'h9cda,
// 16'h9a3a, 16'h99a6, 16'h9b2a, 16'h9eb1,
// 16'ha43c, 16'hab95, 16'hb4b5, 16'hbf49,
// 16'hcb3f, 16'hd836, 16'he608, 16'hf45a,
// 16'h02ec, 16'h116a, 16'h1f96, 16'h2d13,
// 16'h39b1, 16'h451c, 16'h4f25, 16'h5790,
// 16'h5e39, 16'h62f4, 16'h65b2, 16'h665e,
// 16'h64f8, 16'h6186, 16'h5c1a, 16'h54ce,
// 16'h4bd0, 16'h4141, 16'h3568, 16'h2870,
// 16'h1aae, 16'h0c60, 16'hfdcf, 16'hef4d,
// 16'he11f, 16'hd390, 16'hc6ef, 16'hbb6a,
// 16'hb154, 16'ha8d1, 16'ha211, 16'h9d3d,
// 16'h9a63, 16'h999f, 16'h9ae9, 16'h9e43,
// 16'ha395, 16'haac7, 16'hb3b7, 16'hbe2b,
// 16'hc9fe, 16'hd6e1, 16'he49f, 16'hf2e8,
// 16'h0174, 16'h0ffd, 16'h1e2e, 16'h2bc5,
// 16'h387b, 16'h4404, 16'h4e39, 16'h56cc,
// 16'h5da1, 16'h6296, 16'h657f, 16'h6668,
// 16'h6532, 16'h61f6, 16'h5cbb, 16'h559e,
// 16'h4cc8, 16'h425f, 16'h36a4, 16'h29c8,
// 16'h1c16, 16'h0dd2, 16'hff44, 16'hf0bd,
// 16'he285, 16'hd4e2, 16'hc825, 16'hbc83,
// 16'hb245, 16'ha995, 16'ha2ab, 16'h9d9f,
// 16'h9a97, 16'h999b, 16'h9aad, 16'h9dda,
// 16'ha2f2, 16'ha9ff, 16'hb2bc, 16'hbd12,
// 16'hc8bf, 16'hd590, 16'he333, 16'hf17a,
// 16'hfffd, 16'h0e8b, 16'h1cca, 16'h2a71,
// 16'h3742, 16'h42ed, 16'h4d43, 16'h5605,
// 16'h5d08, 16'h622c, 16'h654f, 16'h6665,
// 16'h656c, 16'h625e, 16'h5d57, 16'h566a,
// 16'h4dbb, 16'h437d, 16'h37dc, 16'h2b1c,
// 16'h1d7e, 16'h0f41, 16'h20bc, 16'hf22f,
// 16'he3e8, 16'hd63c, 16'hc959, 16'hbda2,
// 16'hb338, 16'haa61, 16'ha346, 16'h9e0b,
// 16'h9acc, 16'h999b, 16'h9a7e, 16'h9d6c,
// 16'ha25f, 16'ha931, 16'hb1cc, 16'hbbf8,
// 16'hc786, 16'hd43d, 16'he1ce, 16'hf008,
// 16'hfe87, 16'h0d1b, 16'h1b5f, 16'h2921,
// 16'h3602, 16'h41d3, 16'h4c4b, 16'h5537,
// 16'h5c6d, 16'h61bc, 16'h6518, 16'h6661,
// 16'h659b, 16'h62c5, 16'h5dee, 16'h572f,
// 16'h4eae, 16'h4492, 16'h3915, 16'h2c6d,
// 16'h1ee3, 16'h10b2, 16'h0231, 16'hf3a2,
// 16'he550, 16'hd791, 16'hca97, 16'hbec0,
// 16'hb431, 16'hab30, 16'ha3e7, 16'h9e7a,
// 16'h9b08, 16'h99a2, 16'h9a4e, 16'h9d0b,
// 16'ha1c9, 16'ha86e, 16'hb0dd, 16'hbae2,
// 16'hc651, 16'hd2ec, 16'he069, 16'hee99,
// 16'hfd10, 16'h0ba9, 16'h19f9, 16'h27c5,
// 16'h34c7, 16'h40b1, 16'h4b51, 16'h5467,
// 16'h5bc5, 16'h614f, 16'h64d7, 16'h6659,
// 16'h65c7, 16'h6323, 16'h5e82, 16'h57f1,
// 16'h4f99, 16'h45a8, 16'h3a47, 16'h2dc0,
// 16'h2042, 16'h1225, 16'h03a5, 16'hf515,
// 16'he6bb, 16'hd8e6, 16'hcbd9, 16'hbfe2,
// 16'hb52b, 16'hac09, 16'ha486, 16'h9ef4,
// 16'h9b44, 16'h99b1, 16'h9a24, 16'h9cae,
// 16'ha138, 16'ha7b1, 16'hafee, 16'hb9d4,
// 16'hc51c, 16'hd19c, 16'hdf0c, 16'hed23,
// 16'hfba0, 16'h0a33, 16'h188e, 16'h266f,
// 16'h3382, 16'h3f92, 16'h4a4e, 16'h5394,
// 16'h5b1d, 16'h60d7, 16'h6493, 16'h664b,
// 16'h65ee, 16'h637f, 16'h5f0e, 16'h58ad,
// 16'h5084, 16'h46b5, 16'h3b7e, 16'h2f06,
// 16'h21aa, 16'h1390, 16'h051d, 16'hf687,
// 16'he825, 16'hda41, 16'hcd1e, 16'hc102,
// 16'hb633, 16'hacd8, 16'ha539, 16'h9f67,
// 16'h9b8e, 16'h99c1, 16'h9a20, 16'h9c56,
// 16'ha0ad, 16'ha6f5, 16'haf0a, 16'hb8c3,
// 16'hc3ef, 16'hd04e, 16'hddac, 16'hebb4,
// 16'hfa2c, 16'h08be, 16'h1724, 16'h2512,
// 16'h3242, 16'h3e65, 16'h4953, 16'h52b1,
// 16'h5a78, 16'h6056, 16'h644d, 16'h6637,
// 16'h660d, 16'h63d6, 16'h5f96, 16'h5967,
// 16'h5167, 16'h47c3, 16'h3ca9, 16'h3055,
// 16'h2306, 16'h1501, 16'h068f, 16'hf7fd,
// 16'he991, 16'hdb9c, 16'hce64, 16'hc22b,
// 16'hb735, 16'hadb8, 16'ha5e4, 16'h9fe9,
// 16'h9bd8, 16'h99d8, 16'h99e1, 16'h9c03,
// 16'ha027, 16'ha640, 16'hae26, 16'hb7ba,
// 16'hc2c0, 16'hcf07, 16'hdc4b, 16'hea48,
// 16'hf8b6, 16'h074b, 16'h15b6, 16'h23b7,
// 16'h30f7, 16'h3d41, 16'h4846, 16'h51d9,
// 16'h59c1, 16'h5fd9, 16'h63fd, 16'h661e,
// 16'h662a, 16'h6424, 16'h601d, 16'h5a17,
// 16'h524a, 16'h48cb, 16'h3dd4, 16'h319d,
// 16'h2464, 16'h166e, 16'h0804, 16'hf970,
// 16'heaff, 16'hdcfa, 16'hcfac, 16'hc356,
// 16'hb83e, 16'hae97, 16'ha69a, 16'ha06a,
// 16'h9c2b, 16'h99f2, 16'h99c8, 16'h9bb6,
// 16'h9fa4, 16'ha591, 16'had46, 16'hb6b4,
// 16'hc196, 16'hcdc0, 16'hdaef, 16'he8da,
// 16'hf744, 16'h05d3, 16'h144b, 16'h2257,
// 16'h2fae, 16'h3c15, 16'h473a, 16'h50f7,
// 16'h590c, 16'h5f51, 16'h63ad, 16'h65fc,
// 16'h6643, 16'h646f, 16'h609a, 16'h5ac8,
// 16'h5326, 16'h49ce, 16'h3eff, 16'h32e0,
// 16'h25c1, 16'h17db, 16'h0975, 16'hfaea,
// 16'hec69, 16'hde5c, 16'hd0f6, 16'hc483,
// 16'hb94c, 16'haf7c, 16'ha752, 16'ha0f3,
// 16'h9c7f, 16'h9a14, 16'h99b5, 16'h9b6c,
// 16'h9f2a, 16'ha4e1, 16'hac6f, 16'hb5ae,
// 16'hc073, 16'hcc7a, 16'hd993, 16'he771,
// 16'hf5cd, 16'h0461, 16'h12dc, 16'h20f4,
// 16'h2e66, 16'h3ae0, 16'h4631, 16'h500d,
// 16'h5853, 16'h5ec5, 16'h6354, 16'h65db,
// 16'h6651, 16'h64b8, 16'h6111, 16'h5b74,
// 16'h53fc, 16'h4ad3, 16'h401d, 16'h342a,
// 16'h2716, 16'h1947, 16'h0aeb, 16'hfc5a,
// 16'hedde, 16'hdfb9, 16'hd244, 16'hc5b7,
// 16'hba59, 16'hb067, 16'ha80d, 16'ha181,
// 16'h9cdc, 16'h9a38, 16'h99a9, 16'h9b25,
// 16'h9eb6, 16'ha438, 16'hab99, 16'hb4b1,
// 16'hbf4c, 16'hcb3c, 16'hd838, 16'he609,
// 16'hf457, 16'h02ee, 16'h1169, 16'h1f96,
// 16'h2d14, 16'h39b0, 16'h451d, 16'h4f24,
// 16'h5791, 16'h5e37, 16'h62f7, 16'h65af,
// 16'h6662, 16'h64f3, 16'h618a, 16'h5c17,
// 16'h54d1, 16'h4bce, 16'h4143, 16'h3564,
// 16'h2873, 16'h1aae, 16'h0c5e, 16'hfdd3,
// 16'hef48, 16'he122, 16'hd390, 16'hc6ec,
// 16'hbb6e, 16'hb152, 16'ha8d1, 16'ha211,
// 16'h9d3c, 16'h9a66, 16'h999c, 16'h9aec,
// 16'h9e3f, 16'ha398, 16'haac6, 16'hb3b6,
// 16'hbe2e, 16'hc9fb, 16'hd6e4, 16'he49b,
// 16'hf2ea, 16'h0175, 16'h0ffb, 16'h1e31,
// 16'h2bc2, 16'h387c, 16'h4406, 16'h4e36,
// 16'h56ce, 16'h5da1, 16'h6294, 16'h6582,
// 16'h6666, 16'h6533, 16'h61f5, 16'h5cbb,
// 16'h559e, 16'h4cc8, 16'h4260, 16'h36a3,
// 16'h29c9, 16'h1c14, 16'h0dd4, 16'hff42,
// 16'hf0c0, 16'he282, 16'hd4e4, 16'hc825,
// 16'hbc81, 16'hb247, 16'ha994, 16'ha2ac,
// 16'h9d9f, 16'h9a96, 16'h999b, 16'h9ab0,
// 16'h9dd5, 16'ha2f7, 16'ha9fb, 16'hb2be,
// 16'hbd12, 16'hc8be, 16'hd58f, 16'he336,
// 16'hf177, 16'hfffe, 16'h0e8c, 16'h1cc8,
// 16'h2a73, 16'h3742, 16'h42eb, 16'h4d46,
// 16'h5602, 16'h5d0b, 16'h622a, 16'h6550,
// 16'h6666, 16'h6569, 16'h6261, 16'h5d55,
// 16'h566b, 16'h4dbc, 16'h437a, 16'h37df,
// 16'h2b1a, 16'h1d7e, 16'h0f42, 16'h20bc,
// 16'hf22d, 16'he3ec, 16'hd635, 16'hc960,
// 16'hbd9e, 16'hb339, 16'haa62, 16'ha344,
// 16'h9e0c, 16'h9acd, 16'h9999, 16'h9a80,
// 16'h9d6a, 16'ha261, 16'ha92f, 16'hb1ce,
// 16'hbbf7, 16'hc786, 16'hd43d, 16'he1ce,
// 16'hf007, 16'hfe8a, 16'h0d17, 16'h1b63,
// 16'h291d, 16'h3606, 16'h41d1, 16'h4c4b,
// 16'h5538, 16'h5c6a, 16'h61c0, 16'h6515,
// 16'h6663, 16'h659a, 16'h62c6, 16'h5dec,
// 16'h5732, 16'h4eaa, 16'h4496, 16'h3911,
// 16'h2c72, 16'h1ede, 16'h10b6, 16'h022e,
// 16'hf3a3, 16'he551, 16'hd78e, 16'hca9c,
// 16'hbebb, 16'hb434, 16'hab2f, 16'ha3e6,
// 16'h9e7b, 16'h9b08, 16'h99a2, 16'h9a4d,
// 16'h9d0c, 16'ha1c7, 16'ha871, 16'hb0db,
// 16'hbae2, 16'hc652, 16'hd2e9, 16'he06e,
// 16'hee94, 16'hfd14, 16'h0ba6, 16'h19f9,
// 16'h27c7, 16'h34c6, 16'h40b1, 16'h4b50,
// 16'h5468, 16'h5bc5, 16'h614f, 16'h64d6,
// 16'h665a, 16'h65c6, 16'h6326, 16'h5e7e,
// 16'h57f3, 16'h4f9a, 16'h45a5, 16'h3a4c,
// 16'h2dba, 16'h2047, 16'h1221, 16'h03aa,
// 16'hf50f, 16'he6c1, 16'hd8e0, 16'hcbdf,
// 16'hbfdd, 16'hb530, 16'hac03, 16'ha48d,
// 16'h9eed, 16'h9b4a, 16'h99af, 16'h9a23,
// 16'h9cb0, 16'ha136, 16'ha7b2, 16'hafef,
// 16'hb9d2, 16'hc51e, 16'hd19b, 16'hdf0c,
// 16'hed23, 16'hfba0, 16'h0a32, 16'h1890,
// 16'h266c, 16'h3386, 16'h3f8d, 16'h4a53,
// 16'h538f, 16'h5b21, 16'h60d4, 16'h6495,
// 16'h664a, 16'h65ef, 16'h637d, 16'h5f10,
// 16'h58ac, 16'h5084, 16'h46b7, 16'h3b79,
// 16'h2f0d, 16'h21a4, 16'h1394, 16'h051a,
// 16'hf688, 16'he826, 16'hda40, 16'hcd1e,
// 16'hc102, 16'hb632, 16'hacda, 16'ha538,
// 16'h9f66, 16'h9b90, 16'h99bf, 16'h9a01,
// 16'h9c58, 16'ha0a9, 16'ha6f8, 16'haf0a,
// 16'hb8c1, 16'hc3f1, 16'hd04d, 16'hddab,
// 16'hebb7, 16'hfa29, 16'h08bf, 16'h1724,
// 16'h2513, 16'h323e, 16'h3e6c, 16'h494b,
// 16'h52b9, 16'h5a72, 16'h6059, 16'h644d,
// 16'h6635, 16'h6610, 16'h63d3, 16'h5f99,
// 16'h5964, 16'h5169, 16'h47c2, 16'h3caa,
// 16'h3054, 16'h2307, 16'h14ff, 16'h0691,
// 16'hf7fb, 16'he994, 16'hdb99, 16'hce67,
// 16'hc227, 16'hb739, 16'hadb5, 16'ha5e7,
// 16'h9fe6, 16'h9bdb, 16'h99d5, 16'h99e3,
// 16'h9c03, 16'ha026, 16'ha641, 16'hae24,
// 16'hb7bd, 16'hc2bd, 16'hcf0b, 16'hdc47,
// 16'hea4b, 16'hf8b4, 16'h074b, 16'h15b8,
// 16'h23b4, 16'h30fb, 16'h3d3d, 16'h4848,
// 16'h51d9, 16'h59c0, 16'h5fda, 16'h63fc,
// 16'h661f, 16'h6629, 16'h6427, 16'h6018,
// 16'h5a1c, 16'h5247, 16'h48cc, 16'h3dd4,
// 16'h319d, 16'h2464, 16'h166e, 16'h0804,
// 16'hf971, 16'heafe, 16'hdcfa, 16'hcfac,
// 16'hc355, 16'hb841, 16'hae94, 16'ha69d,
// 16'ha067, 16'h9c2c, 16'h99f3, 16'h99c6,
// 16'h9bb9, 16'h9fa2, 16'ha591, 16'had47,
// 16'hb6b3, 16'hc196, 16'hcdc2, 16'hdaeb,
// 16'he8df, 16'hf740, 16'h05d5, 16'h144c,
// 16'h2253, 16'h2fb3, 16'h3c11, 16'h473d,
// 16'h50f5, 16'h590e, 16'h5f4e, 16'h63af,
// 16'h65fc, 16'h6642, 16'h6470, 16'h609a,
// 16'h5ac7, 16'h5327, 16'h49ce, 16'h3efd,
// 16'h32e3, 16'h25bf, 16'h17dc, 16'h0975,
// 16'hfae9, 16'hec6a, 16'hde5c, 16'hd0f4,
// 16'hc487, 16'hb948, 16'haf7f, 16'ha750,
// 16'ha0f3, 16'h9c81, 16'h9a12, 16'h99b6,
// 16'h9b6c, 16'h9f29, 16'ha4e3, 16'hac6d,
// 16'hb5b0, 16'hc071, 16'hcc7b, 16'hd993,
// 16'he772, 16'hf5cc, 16'h0461, 16'h12dc,
// 16'h20f4, 16'h2e66, 16'h3ae1, 16'h462f,
// 16'h500f, 16'h5851, 16'h5ec7, 16'h6353,
// 16'h65da, 16'h6653, 16'h64b6, 16'h6113,
// 16'h5b73, 16'h53fc, 16'h4ad2, 16'h4020,
// 16'h3427, 16'h2718, 16'h1946, 16'h0aeb,
// 16'hfc5b, 16'heddc, 16'hdfbb, 16'hd243,
// 16'hc5b7, 16'hba5a, 16'hb065, 16'ha80f,
// 16'ha180, 16'h9cdc, 16'h9a39, 16'h99a6,
// 16'h9b2a, 16'h9eb1, 16'ha43c, 16'hab97,
// 16'hb4b1, 16'hbf4d, 16'hcb3b, 16'hd838,
// 16'he609, 16'hf458, 16'h02ee, 16'h1169,
// 16'h1f95, 16'h2d14, 16'h39b1, 16'h451c,
// 16'h4f25, 16'h5790, 16'h5e39, 16'h62f3,
// 16'h65b5, 16'h665a, 16'h64fc, 16'h6183,
// 16'h5c1a, 16'h54d2, 16'h4bca, 16'h4147,
// 16'h3563, 16'h2872, 16'h1aaf, 16'h0c5e,
// 16'hfdd0, 16'hef4d, 16'he11e, 16'hd392,
// 16'hc6ec, 16'hbb6d, 16'hb152, 16'ha8d2,
// 16'ha211, 16'h9d3b, 16'h9a67, 16'h999b,
// 16'h9aec, 16'h9e41, 16'ha395, 16'haac9,
// 16'hb3b4, 16'hbe2e, 16'hc9fc, 16'hd6e2,
// 16'he49f, 16'hf2e6, 16'h0178, 16'h0ff9,
// 16'h1e31, 16'h2bc3, 16'h387c, 16'h4405,
// 16'h4e38, 16'h56cb, 16'h5da3, 16'h6294,
// 16'h6581, 16'h6667, 16'h6532, 16'h61f6,
// 16'h5cba, 16'h55a0, 16'h4cc6, 16'h4262,
// 16'h36a1, 16'h29c9, 16'h1c16, 16'h0dd2,
// 16'hff44, 16'hf0be, 16'he282, 16'hd4e6,
// 16'hc821, 16'hbc86, 16'hb242, 16'ha998,
// 16'ha2a9, 16'h9da0, 16'h9a98, 16'h9996,
// 16'h9ab5, 16'h9dd2, 16'ha2f9, 16'ha9fa,
// 16'hb2bd, 16'hbd14, 16'hc8bc, 16'hd593,
// 16'he331, 16'hf17a, 16'hfffe, 16'h0e8a,
// 16'h1ccb, 16'h2a70, 16'h3743, 16'h42ec,
// 16'h4d45, 16'h5602, 16'h5d0b, 16'h622b,
// 16'h654e, 16'h6669, 16'h6566, 16'h6263,
// 16'h5d54, 16'h566c, 16'h4dba, 16'h437d,
// 16'h37dc, 16'h2b1c, 16'h1d7e, 16'h0f40,
// 16'h20be, 16'hf22c, 16'he3ec, 16'hd637,
// 16'hc95d, 16'hbda0, 16'hb339, 16'haa5f,
// 16'ha349, 16'h9e07, 16'h9ad0, 16'h9999,
// 16'h9a7d, 16'h9d6e, 16'ha25c, 16'ha935,
// 16'hb1c8, 16'hbbfb, 16'hc784, 16'hd43e,
// 16'he1ce, 16'hf007, 16'hfe88, 16'h0d1b,
// 16'h1b5f, 16'h2922, 16'h3620, 16'h41d4,
// 16'h4c4b, 16'h5538, 16'h5c6b, 16'h61be,
// 16'h6515, 16'h6664, 16'h659a, 16'h62c5,
// 16'h5dee, 16'h572e, 16'h4eaf, 16'h4491,
// 16'h3917, 16'h2c6c, 16'h1ee2, 16'h10b4,
// 16'h022f, 16'hf3a3, 16'he551, 16'hd78e,
// 16'hca9b, 16'hbebc, 16'hb434, 16'hab2f,
// 16'ha3e7, 16'h9e79, 16'h9b08, 16'h99a3,
// 16'h9a4e, 16'h9d0b, 16'ha1c9, 16'ha86c,
// 16'hb0e0, 16'hbade, 16'hc657, 16'hd2e4,
// 16'he073, 16'hee8f, 16'hfd18, 16'h0ba3,
// 16'h19fc, 16'h27c5, 16'h34c8, 16'h40af,
// 16'h4b52, 16'h5466, 16'h5bc8, 16'h614c,
// 16'h64d9, 16'h6657, 16'h65c9, 16'h6323,
// 16'h5e81, 16'h57f1, 16'h4f9a, 16'h45a6,
// 16'h3a4b, 16'h2dbb, 16'h2047, 16'h1221,
// 16'h03a8, 16'hf513, 16'he6bc, 16'hd8e6,
// 16'hcbda, 16'hbfdf, 16'hb531, 16'hac01,
// 16'ha48e, 16'h9eed, 16'h9b4a, 16'h99ad,
// 16'h9a27, 16'h9cab, 16'ha13b, 16'ha7ad,
// 16'haff4, 16'hb9cd, 16'hc522, 16'hd199,
// 16'hdf0c, 16'hed24, 16'hfba0, 16'h0a31,
// 16'h1892, 16'h266a, 16'h3387, 16'h3f8e,
// 16'h4a50, 16'h5393, 16'h5b1d, 16'h60d7,
// 16'h6495, 16'h6649, 16'h65ee, 16'h637f,
// 16'h5f0e, 16'h58ae, 16'h5084, 16'h46b5,
// 16'h3b7c, 16'h2f09, 16'h21a7, 16'h1392,
// 16'h051c, 16'hf686, 16'he829, 16'hda3c,
// 16'hcd21, 16'hc101, 16'hb632, 16'hacda,
// 16'ha538, 16'h9f66, 16'h9b91, 16'h99be,
// 16'h9a01, 16'h9c56, 16'ha0ad, 16'ha6f5,
// 16'haf0b, 16'hb8c1, 16'hc3f1, 16'hd04d,
// 16'hddac, 16'hebb5, 16'hfa2a, 16'h08c0,
// 16'h1723, 16'h2513, 16'h3240, 16'h3e68,
// 16'h494e, 16'h52b7, 16'h5a73, 16'h605a,
// 16'h644b, 16'h6637, 16'h660e, 16'h63d6,
// 16'h5f95, 16'h5967, 16'h5168, 16'h47c3,
// 16'h3ca8, 16'h3057, 16'h2302, 16'h1505,
// 16'h068c, 16'hf7ff, 16'he990, 16'hdb9c,
// 16'hce65, 16'hc228, 16'hb739, 16'hadb4,
// 16'ha5e8, 16'h9fe6, 16'h9bd9, 16'h99d7,
// 16'h99e2, 16'h9c03, 16'ha027, 16'ha63e,
// 16'hae29, 16'hb7b7, 16'hc2c2, 16'hcf07,
// 16'hdc4a, 16'hea49, 16'hf8b6, 16'h074a,
// 16'h15b7, 16'h23b7, 16'h30f7, 16'h3d41,
// 16'h4847, 16'h51d7, 16'h59c4, 16'h5fd5,
// 16'h6401, 16'h661c, 16'h662a, 16'h6426,
// 16'h6019, 16'h5a1b, 16'h5248, 16'h48cc,
// 16'h3dd2, 16'h31a0, 16'h2461, 16'h1671,
// 16'h0801, 16'hf973, 16'heafd, 16'hdcfc,
// 16'hcfa9, 16'hc358, 16'hb83e, 16'hae97,
// 16'ha69b, 16'ha068, 16'h9c2c, 16'h99f2,
// 16'h99c8, 16'h9bb6, 16'h9fa5, 16'ha58f,
// 16'had48, 16'hb6b2, 16'hc197, 16'hcdc0,
// 16'hdaef, 16'he8db, 16'hf741, 16'h05d7,
// 16'h1447, 16'h225b, 16'h2fab, 16'h3c17,
// 16'h4739, 16'h50f8, 16'h590b, 16'h5f52,
// 16'h63ab, 16'h65ff, 16'h6640, 16'h6472,
// 16'h6098, 16'h5ac8, 16'h5326, 16'h49cf,
// 16'h3efd, 16'h32e3, 16'h25bf, 16'h17da,
// 16'h0979, 16'hfae4, 16'hec6f, 16'hde58,
// 16'hd0f7, 16'hc485, 16'hb949, 16'haf7e,
// 16'ha750, 16'ha0f5, 16'h9c7e, 16'h9a15,
// 16'h99b3, 16'h9b6e, 16'h9f29, 16'ha4e2,
// 16'hac6e, 16'hb5af, 16'hc072, 16'hcc7a,
// 16'hd994, 16'he771, 16'hf5cc, 16'h0462,
// 16'h12da, 16'h20f6, 16'h2e65, 16'h3ae1,
// 16'h4630, 16'h500e, 16'h5851, 16'h5ec8,
// 16'h6351, 16'h65dc, 16'h6652, 16'h64b7,
// 16'h6112, 16'h5b73, 16'h53fc, 16'h4ad2,
// 16'h4021, 16'h3425, 16'h271a, 16'h1945,
// 16'h0aec, 16'hfc5a, 16'heddd, 16'hdfba,
// 16'hd245, 16'hc5b5, 16'hba5b, 16'hb065,
// 16'ha80f, 16'ha181, 16'h9cd9, 16'h9a3d,
// 16'h99a2, 16'h9b2d, 16'h9eb0, 16'ha43b,
// 16'hab98, 16'hb4b1, 16'hbf4d, 16'hcb3a,
// 16'hd83a, 16'he607, 16'hf459, 16'h02ee,
// 16'h1167, 16'h1f99, 16'h2d11, 16'h39b2,
// 16'h451c, 16'h4f23, 16'h5794, 16'h5e35,
// 16'h62f7, 16'h65b1, 16'h665d, 16'h64fa,
// 16'h6184, 16'h5c1b, 16'h54cf, 16'h4bce,
// 16'h4144, 16'h3563, 16'h2875, 16'h1aaa,
// 16'h0c63, 16'hfdcc, 16'hef50, 16'he11c,
// 16'hd393, 16'hc6eb, 16'hbb6e, 16'hb152,
// 16'ha8d2, 16'ha211, 16'h9d3b, 16'h9a67,
// 16'h999b, 16'h9aec, 16'h9e41, 16'ha395,
// 16'haac9, 16'hb3b4, 16'hbe2e, 16'hc9fc,
// 16'hd6e2, 16'he49f, 16'hf2e6, 16'h0177,
// 16'h0ffb, 16'h1e2f, 16'h2bc6, 16'h3879,
// 16'h4406, 16'h4e37, 16'h56cd, 16'h5da2,
// 16'h6294, 16'h6581, 16'h6666, 16'h6534,
// 16'h61f4, 16'h5cbc, 16'h559d, 16'h4cc9,
// 16'h425f, 16'h36a4, 16'h29c8, 16'h1c15,
// 16'h0dd2, 16'hff46, 16'hf0bc, 16'he284,
// 16'hd4e4, 16'hc822, 16'hbc87, 16'hb241,
// 16'ha999, 16'ha2a7, 16'h9da3, 16'h9a94,
// 16'h999b, 16'h9ab0, 16'h9dd6, 16'ha2f6,
// 16'ha9fb, 16'hb2bf, 16'hbd0f, 16'hc8c3,
// 16'hd58a, 16'he33a, 16'hf173, 16'h2002,
// 16'h0e88, 16'h1ccc, 16'h2a70, 16'h3743,
// 16'h42eb, 16'h4d45, 16'h5603, 16'h5d0b,
// 16'h622a, 16'h6550, 16'h6665, 16'h656b,
// 16'h625f, 16'h5d57, 16'h5669, 16'h4dbd,
// 16'h437a, 16'h37df, 16'h2b1a, 16'h1d7e,
// 16'h0f42, 16'h20bc, 16'hf22d, 16'he3ec,
// 16'hd636, 16'hc95f, 16'hbd9e, 16'hb339,
// 16'haa63, 16'ha343, 16'h9e0d, 16'h9acb,
// 16'h999b, 16'h9a7f, 16'h9d6a, 16'ha261,
// 16'ha930, 16'hb1cc, 16'hbbf9, 16'hc785,
// 16'hd43c, 16'he1d1, 16'hf004, 16'hfe8b,
// 16'h0d18, 16'h1b62, 16'h291d, 16'h3606,
// 16'h41d0, 16'h4c4d, 16'h5537, 16'h5c6a,
// 16'h61c0, 16'h6515, 16'h6663, 16'h659a,
// 16'h62c5, 16'h5dee, 16'h572f, 16'h4eae,
// 16'h4491, 16'h3917, 16'h2c6c, 16'h1ee3,
// 16'h10b1, 16'h0233, 16'hf39f, 16'he554,
// 16'hd78d, 16'hca9a, 16'hbebe, 16'hb432,
// 16'hab30, 16'ha3e7, 16'h9e7a, 16'h9b06,
// 16'h99a5, 16'h9a4c, 16'h9d0c, 16'ha1c9,
// 16'ha86d, 16'hb0de, 16'hbae2, 16'hc650,
// 16'hd2eb, 16'he06d, 16'hee94, 16'hfd15,
// 16'h0ba5, 16'h19fb, 16'h27c3, 16'h34ca,
// 16'h40af, 16'h4b52, 16'h5465, 16'h5bc9,
// 16'h614b, 16'h64d8, 16'h665b, 16'h65c3,
// 16'h6329, 16'h5e7d, 16'h57f2, 16'h4f9a,
// 16'h45a7, 16'h3a48, 16'h2dbf, 16'h2043,
// 16'h1224, 16'h03a6, 16'hf514, 16'he6bc,
// 16'hd8e5, 16'hcbdb, 16'hbfdf, 16'hb52f,
// 16'hac05, 16'ha48a, 16'h9eef, 16'h9b4a,
// 16'h99ad, 16'h9a26, 16'h9cad, 16'ha138,
// 16'ha7b1, 16'haff0, 16'hb9d2, 16'hc51d,
// 16'hd19c, 16'hdf0b, 16'hed24, 16'hfba0,
// 16'h0a32, 16'h1890, 16'h266c, 16'h3386,
// 16'h3f8d, 16'h4a52, 16'h5392, 16'h5b1d,
// 16'h60d8, 16'h6493, 16'h664a, 16'h65ef,
// 16'h637d, 16'h5f0f, 16'h58ae, 16'h5083,
// 16'h46b7, 16'h3b7a, 16'h2f0b, 16'h21a4,
// 16'h1396, 16'h0517, 16'hf68d, 16'he820,
// 16'hda46, 16'hcd18, 16'hc108, 16'hb62d,
// 16'hacdd, 16'ha536, 16'h9f68, 16'h9b8f,
// 16'h99bf, 16'h9a01, 16'h9c56, 16'ha0ac,
// 16'ha6f7, 16'haf08, 16'hb8c4, 16'hc3ee,
// 16'hd04f, 16'hddab, 16'hebb5, 16'hfa2b,
// 16'h08be, 16'h1725, 16'h2511, 16'h3241,
// 16'h3e68, 16'h494f, 16'h52b6, 16'h5a73,
// 16'h605a, 16'h644b, 16'h6637, 16'h660f,
// 16'h63d4, 16'h5f97, 16'h5966, 16'h5168,
// 16'h47c2, 16'h3caa, 16'h3054, 16'h2307,
// 16'h14ff, 16'h0692, 16'hf7f9, 16'he995,
// 16'hdb99, 16'hce66, 16'hc229, 16'hb737,
// 16'hadb7, 16'ha5e4, 16'h9fe9, 16'h9bd8,
// 16'h99d8, 16'h99e1, 16'h9c03, 16'ha027,
// 16'ha63f, 16'hae27, 16'hb7ba, 16'hc2bf,
// 16'hcf09, 16'hdc49, 16'hea49, 16'hf8b6,
// 16'h074a, 16'h15b8, 16'h23b4, 16'h30fb,
// 16'h3d3d, 16'h4849, 16'h51d8, 16'h59c1,
// 16'h5fd9, 16'h63fc, 16'h6620, 16'h6628,
// 16'h6428, 16'h6017, 16'h5a1d, 16'h5246,
// 16'h48cd, 16'h3dd3, 16'h319d, 16'h2465,
// 16'h166d, 16'h0804, 16'hf972, 16'heafc,
// 16'hdcfd, 16'hcfa9, 16'hc358, 16'hb83d,
// 16'hae98, 16'ha69a, 16'ha069, 16'h9c2c,
// 16'h99f1, 16'h99c9, 16'h9bb5, 16'h9fa6,
// 16'ha58d, 16'had4b, 16'hb6b0, 16'hc198,
// 16'hcdc0, 16'hdaed, 16'he8dd, 16'hf741,
// 16'h05d6, 16'h1449, 16'h2258, 16'h2fae,
// 16'h3c13, 16'h473e, 16'h50f4, 16'h590e,
// 16'h5f4f, 16'h63ad, 16'h65fe, 16'h6641,
// 16'h6471, 16'h6098, 16'h5ac9, 16'h5326,
// 16'h49ce, 16'h3efe, 16'h32e1, 16'h25c2,
// 16'h17d8, 16'h097a, 16'hfae4, 16'hec6d,
// 16'hde5b, 16'hd0f4, 16'hc488, 16'hb947,
// 16'haf80, 16'ha74e, 16'ha0f6, 16'h9c7e,
// 16'h9a14, 16'h99b6, 16'h9b6a, 16'h9f2c,
// 16'ha4e0, 16'hac6f, 16'hb5af, 16'hc071,
// 16'hcc7b, 16'hd995, 16'he76e, 16'hf5d0,
// 16'h045e, 16'h12de, 16'h20f3, 16'h2e67,
// 16'h3adf, 16'h4632, 16'h500c, 16'h5853,
// 16'h5ec6, 16'h6354, 16'h65d9, 16'h6654,
// 16'h64b5, 16'h6114, 16'h5b71, 16'h5420,
// 16'h4acc, 16'h4027, 16'h341f, 16'h2720,
// 16'h193f, 16'h0af0, 16'hfc59, 16'heddb,
// 16'hdfbe, 16'hd240, 16'hc5b9, 16'hba58,
// 16'hb067, 16'ha80e, 16'ha181, 16'h9cda,
// 16'h9a3b, 16'h99a5, 16'h9b29, 16'h9eb3,
// 16'ha43a, 16'hab98, 16'hb4b1, 16'hbf4c,
// 16'hcb3c, 16'hd838, 16'he609, 16'hf458,
// 16'h02ec, 16'h116c, 16'h1f92, 16'h2d18,
// 16'h39ad, 16'h451e, 16'h4f23, 16'h5792,
// 16'h5e38, 16'h62f4, 16'h65b2, 16'h665e,
// 16'h64f8, 16'h6187, 16'h5c17, 16'h54d3,
// 16'h4bcb, 16'h4145, 16'h3564, 16'h2872,
// 16'h1ab0, 16'h0c5d, 16'hfdd0, 16'hef4d,
// 16'he11d, 16'hd394, 16'hc6eb, 16'hbb6c,
// 16'hb156, 16'ha8cc, 16'ha216, 16'h9d39,
// 16'h9a66, 16'h999e, 16'h9ae9, 16'h9e42,
// 16'ha397, 16'haac5, 16'hb3b7, 16'hbe2d,
// 16'hc9fc, 16'hd6e3, 16'he49c, 16'hf2ea,
// 16'h0173, 16'h0ffe, 16'h1e2d, 16'h2bc7,
// 16'h3878, 16'h4408, 16'h4e35, 16'h56cd,
// 16'h5da4, 16'h6291, 16'h6585, 16'h6662,
// 16'h6536, 16'h61f4, 16'h5cbb, 16'h559f,
// 16'h4cc6, 16'h4262, 16'h36a2, 16'h29c9,
// 16'h1c15, 16'h0dd2, 16'hff44, 16'hf0bf,
// 16'he282, 16'hd4e5, 16'hc822, 16'hbc85,
// 16'hb243, 16'ha998, 16'ha2a8, 16'h9da1,
// 16'h9a96, 16'h999a, 16'h9ab0, 16'h9dd7,
// 16'ha2f3, 16'ha9ff, 16'hb2bb, 16'hbd14,
// 16'hc8be, 16'hd58e, 16'he336, 16'hf177,
// 16'hffff, 16'h0e8c, 16'h1cc6, 16'h2a76,
// 16'h373e, 16'h42ef, 16'h4d43, 16'h5603,
// 16'h5d0a, 16'h622c, 16'h654e, 16'h6667,
// 16'h6569, 16'h625f, 16'h5d59, 16'h5667,
// 16'h4dbf, 16'h4378, 16'h37df, 16'h2b1c,
// 16'h1d7c, 16'h0f44, 16'h20b9, 16'hf230,
// 16'he3ea, 16'hd637, 16'hc95e, 16'hbd9f,
// 16'hb339, 16'haa62, 16'ha344, 16'h9e0c,
// 16'h9acb, 16'h999d, 16'h9a7b, 16'h9d70,
// 16'ha25a, 16'ha936, 16'hb1c9, 16'hbbf7,
// 16'hc78b, 16'hd436, 16'he1d5, 16'hf002,
// 16'hfe8b, 16'h0d19, 16'h1b61, 16'h291f,
// 16'h3602, 16'h41d5, 16'h4c48, 16'h553b,
// 16'h5c69, 16'h61be, 16'h6517, 16'h6662,
// 16'h659b, 16'h62c5, 16'h5dec, 16'h5731,
// 16'h4ead, 16'h4492, 16'h3917, 16'h2c6a,
// 16'h1ee4, 16'h10b3, 16'h0230, 16'hf3a2,
// 16'he551, 16'hd78f, 16'hca99, 16'hbec0,
// 16'hb42f, 16'hab33, 16'ha3e3, 16'h9e7d,
// 16'h9b06, 16'h99a4, 16'h9a4c, 16'h9d0d,
// 16'ha1c7, 16'ha86f, 16'hb0dc, 16'hbae3,
// 16'hc651, 16'hd2ea, 16'he06e, 16'hee92,
// 16'hfd17, 16'h0ba4, 16'h19fa, 16'h27c7,
// 16'h34c5, 16'h40b3, 16'h4b4f, 16'h5468,
// 16'h5bc6, 16'h614e, 16'h64d7, 16'h6659,
// 16'h65c8, 16'h6323, 16'h5e82, 16'h57ef,
// 16'h4f9c, 16'h45a6, 16'h3a48, 16'h2dc0,
// 16'h2040, 16'h1229, 16'h03a2, 16'hf515,
// 16'he6bc, 16'hd8e5, 16'hcbdc, 16'hbfde,
// 16'hb52f, 16'hac04, 16'ha48c, 16'h9eef,
// 16'h9b49, 16'h99ac, 16'h9a28, 16'h9cab,
// 16'ha13b, 16'ha7ae, 16'haff2, 16'hb9ce,
// 16'hc522, 16'hd198, 16'hdf0f, 16'hed21,
// 16'hfba1, 16'h0a31, 16'h1891, 16'h266c,
// 16'h3385, 16'h3f8f, 16'h4a51, 16'h5391,
// 16'h5b1f, 16'h60d5, 16'h6495, 16'h664b,
// 16'h65ec, 16'h6381, 16'h5f0c, 16'h58af,
// 16'h5083, 16'h46b7, 16'h3b79, 16'h2f0c,
// 16'h21a5, 16'h1393, 16'h051c, 16'hf686,
// 16'he826, 16'hda41, 16'hcd1d, 16'hc104,
// 16'hb630, 16'hacdb, 16'ha536, 16'h9f6a,
// 16'h9b8d, 16'h99c1, 16'h99ff, 16'h9c57,
// 16'ha0ac, 16'ha6f7, 16'haf08, 16'hb8c5,
// 16'hc3eb, 16'hd053, 16'hdda7, 16'hebb9,
// 16'hfa28, 16'h08c0, 16'h1723, 16'h2512,
// 16'h3242, 16'h3e66, 16'h4950, 16'h52b6,
// 16'h5a72, 16'h605b, 16'h644a, 16'h6639,
// 16'h660b, 16'h63d9, 16'h5f91, 16'h596d,
// 16'h5162, 16'h47c7, 16'h3ca6, 16'h3057,
// 16'h2304, 16'h1503, 16'h068e, 16'hf7fd,
// 16'he992, 16'hdb9b, 16'hce63, 16'hc22d,
// 16'hb734, 16'hadb8, 16'ha5e5, 16'h9fe7,
// 16'h9bd9, 16'h99d8, 16'h99e1, 16'h9c02,
// 16'ha02a, 16'ha63b, 16'hae2c, 16'hb7b4,
// 16'hc2c5, 16'hcf04, 16'hdc4c, 16'hea49,
// 16'hf8b4, 16'h074c, 16'h15b6, 16'h23b6,
// 16'h30f9, 16'h3d3f, 16'h4847, 16'h51d9,
// 16'h59c1, 16'h5fd9, 16'h63fd, 16'h661d,
// 16'h662b, 16'h6425, 16'h601b, 16'h5a19,
// 16'h5248, 16'h48cd, 16'h3dd1, 16'h31a1,
// 16'h2461, 16'h166e, 16'h0807, 16'hf96c,
// 16'heb04, 16'hdcf5, 16'hcfaf, 16'hc354,
// 16'hb840, 16'hae96, 16'ha69c, 16'ha067,
// 16'h9c2c, 16'h99f2, 16'h99c9, 16'h9bb5,
// 16'h9fa6, 16'ha58c, 16'had4c, 16'hb6af,
// 16'hc19a, 16'hcdbd, 16'hdaf0, 16'he8da,
// 16'hf744, 16'h05d3, 16'h144c, 16'h2255,
// 16'h2faf, 16'h3c15, 16'h473a, 16'h50f8,
// 16'h590b, 16'h5f51, 16'h63ac, 16'h65fe,
// 16'h6640, 16'h6474, 16'h6094, 16'h5acd,
// 16'h5322, 16'h49d1, 16'h3efc, 16'h32e3,
// 16'h25c0, 16'h17d9, 16'h097a, 16'hfae3,
// 16'hec6f, 16'hde5a, 16'hd0f4, 16'hc487,
// 16'hb949, 16'haf7c, 16'ha754, 16'ha0f0,
// 16'h9c82, 16'h9a12, 16'h99b6, 16'h9b6c,
// 16'h9f2a, 16'ha4e0, 16'hac71, 16'hb5ad,
// 16'hc073, 16'hcc7a, 16'hd993, 16'he772,
// 16'hf5cc, 16'h0461, 16'h12dc, 16'h20f5,
// 16'h2e64, 16'h3ae2, 16'h462f, 16'h5010,
// 16'h5850, 16'h5ec8, 16'h6351, 16'h65dc,
// 16'h6652, 16'h64b7, 16'h6112, 16'h5b74,
// 16'h53fb, 16'h4ad3, 16'h401e, 16'h3428,
// 16'h2719, 16'h1946, 16'h0ae9, 16'hfc5e,
// 16'hedd8, 16'hdfc0, 16'hd23f, 16'hc5ba,
// 16'hba57, 16'hb068, 16'ha80d, 16'ha182,
// 16'h9cd9, 16'h9a3b, 16'h99a6, 16'h9b28,
// 16'h9eb5, 16'ha437, 16'hab9a, 16'hb4b0,
// 16'hbf4e, 16'hcb3a, 16'hd839, 16'he607,
// 16'hf45b, 16'h02ea, 16'h116e, 16'h1f90,
// 16'h2d18, 16'h39af, 16'h451c, 16'h4f25,
// 16'h5791, 16'h5e38, 16'h62f4, 16'h65b3,
// 16'h665c, 16'h64fb, 16'h6183, 16'h5c1b,
// 16'h54d0, 16'h4bcd, 16'h4144, 16'h3565,
// 16'h2871, 16'h1aaf, 16'h0c60, 16'hfdcd,
// 16'hef50, 16'he11b, 16'hd395, 16'hc6e9,
// 16'hbb6f, 16'hb153, 16'ha8ce, 16'ha216,
// 16'h9d37, 16'h9a69, 16'h999b, 16'h9aeb,
// 16'h9e42, 16'ha394, 16'haac9, 16'hb3b5,
// 16'hbe2d, 16'hc9fd, 16'hd6e1, 16'he49f,
// 16'hf2e7, 16'h0177, 16'h0ffa, 16'h1e2f,
// 16'h2bc6, 16'h3878, 16'h440a, 16'h4e32,
// 16'h56d0, 16'h5da0, 16'h6296, 16'h657f,
// 16'h6669, 16'h6530, 16'h61f7, 16'h5cbb,
// 16'h559e, 16'h4cc7, 16'h4262, 16'h36a0,
// 16'h29cb, 16'h1c14, 16'h0dd2, 16'hff46,
// 16'hf0bb, 16'he285, 16'hd4e3, 16'hc824,
// 16'hbc83, 16'hb246, 16'ha993, 16'ha2ad,
// 16'h9d9f, 16'h9a96, 16'h999b, 16'h9aaf,
// 16'h9dd6, 16'ha2f7, 16'ha9fa, 16'hb2c0,
// 16'hbd10, 16'hc8c0, 16'hd58e, 16'he335,
// 16'hf178, 16'hffff, 16'h0e8a, 16'h1cca,
// 16'h2a72, 16'h3741, 16'h42ed, 16'h4d44,
// 16'h5602, 16'h5d0c, 16'h622a, 16'h654f,
// 16'h6667, 16'h6569, 16'h625f, 16'h5d58,
// 16'h5668, 16'h4dbe, 16'h437a, 16'h37de,
// 16'h2b1c, 16'h1d7b, 16'h0f45, 16'h20b9,
// 16'hf230, 16'he3e9, 16'hd639, 16'hc95c,
// 16'hbda1, 16'hb337, 16'haa62, 16'ha346,
// 16'h9e0a, 16'h9acd, 16'h999a, 16'h9a7e,
// 16'h9d6d, 16'ha25d, 16'ha933, 16'hb1cb,
// 16'hbbf8, 16'hc787, 16'hd43b, 16'he1d0,
// 16'hf006, 16'hfe8a, 16'h0d18, 16'h1b62,
// 16'h291e, 16'h3603, 16'h41d4, 16'h4c4a,
// 16'h5538, 16'h5c6b, 16'h61be, 16'h6516,
// 16'h6663, 16'h659a, 16'h62c6, 16'h5dec,
// 16'h5731, 16'h4eac, 16'h4494, 16'h3915,
// 16'h2c6b, 16'h1ee4, 16'h10b2, 16'h0231,
// 16'hf3a2, 16'he550, 16'hd78f, 16'hca9b,
// 16'hbebb, 16'hb436, 16'hab2c, 16'ha3e9,
// 16'h9e7a, 16'h9b06, 16'h99a4, 16'h9a4d,
// 16'h9d0b, 16'ha1ca, 16'ha86d, 16'hb0dc,
// 16'hbae4, 16'hc64f, 16'hd2ed, 16'he06a,
// 16'hee96, 16'hfd14, 16'h0ba5, 16'h19fb,
// 16'h27c5, 16'h34c6, 16'h40b3, 16'h4b4f,
// 16'h5467, 16'h5bc8, 16'h614b, 16'h64da,
// 16'h6657, 16'h65c8, 16'h6324, 16'h5e81,
// 16'h57f0, 16'h4f9c, 16'h45a4, 16'h3a4c,
// 16'h2dbb, 16'h2046, 16'h1222, 16'h03a8,
// 16'hf513, 16'he6bb, 16'hd8e8, 16'hcbd6,
// 16'hbfe5, 16'hb52a, 16'hac07, 16'ha48a,
// 16'h9eef, 16'h9b4a, 16'h99ac, 16'h9a27,
// 16'h9cac, 16'ha13a, 16'ha7af, 16'haff0,
// 16'hb9d3, 16'hc51b, 16'hd19f, 16'hdf09,
// 16'hed24, 16'hfba1, 16'h0a30, 16'h1891,
// 16'h266e, 16'h3382, 16'h3f91, 16'h4a50,
// 16'h5391, 16'h5b20, 16'h60d4, 16'h6496,
// 16'h6649, 16'h65ef, 16'h637e, 16'h5f0e,
// 16'h58ae, 16'h5082, 16'h46b9, 16'h3b78,
// 16'h2f0d, 16'h21a3, 16'h1395, 16'h051a,
// 16'hf689, 16'he824, 16'hda41, 16'hcd1e,
// 16'hc103, 16'hb632, 16'hacd8, 16'ha53a,
// 16'h9f64, 16'h9b94, 16'h99bb, 16'h9a05,
// 16'h9c52, 16'ha0af, 16'ha6f4, 16'haf0c,
// 16'hb8c1, 16'hc3f0, 16'hd04d, 16'hddac,
// 16'hebb5, 16'hfa2c, 16'h08bd, 16'h1724,
// 16'h2514, 16'h323d, 16'h3e6d, 16'h4949,
// 16'h52bc, 16'h5a6f, 16'h605b, 16'h644c,
// 16'h6635, 16'h6610, 16'h63d5, 16'h5f95,
// 16'h5968, 16'h5166, 16'h47c4, 16'h3ca9,
// 16'h3055, 16'h2306, 16'h1520, 16'h0691,
// 16'hf7fb, 16'he992, 16'hdb9d, 16'hce62,
// 16'hc22e, 16'hb731, 16'hadbb, 16'ha5e3,
// 16'h9fe9, 16'h9bd9, 16'h99d6, 16'h99e2,
// 16'h9c03, 16'ha027, 16'ha63f, 16'hae28,
// 16'hb7b8, 16'hc2c1, 16'hcf06, 16'hdc4c,
// 16'hea47, 16'hf8b8, 16'h0748, 16'h15b8,
// 16'h23b6, 16'h30f8, 16'h3d41, 16'h4846,
// 16'h51d8, 16'h59c2, 16'h5fd8, 16'h63ff,
// 16'h661c, 16'h662b, 16'h6424, 16'h601d,
// 16'h5a17, 16'h524b, 16'h48c9, 16'h3dd5,
// 16'h319e, 16'h2463, 16'h166e, 16'h0805,
// 16'hf96e, 16'heb02, 16'hdcf8, 16'hcfac,
// 16'hc357, 16'hb83d, 16'hae97, 16'ha69d,
// 16'ha065, 16'h9c30, 16'h99ee, 16'h99cb,
// 16'h9bb4, 16'h9fa6, 16'ha58e, 16'had49,
// 16'hb6b2, 16'hc196, 16'hcdc2, 16'hdaec,
// 16'he8dd, 16'hf742, 16'h05d3, 16'h144d,
// 16'h2254, 16'h2fb1, 16'h3c12, 16'h473e,
// 16'h50f3, 16'h590f, 16'h5f4f, 16'h63ad,
// 16'h65fe, 16'h6641, 16'h6471, 16'h6098,
// 16'h5ac9, 16'h5325, 16'h49d0, 16'h3efc,
// 16'h32e3, 16'h25bf, 16'h17da, 16'h0979,
// 16'hfae5, 16'hec6c, 16'hde5c, 16'hd0f2,
// 16'hc48a, 16'hb946, 16'haf7f, 16'ha751,
// 16'ha0f2, 16'h9c81, 16'h9a13, 16'h99b5,
// 16'h9b6c, 16'h9f2a, 16'ha4e1, 16'hac6f,
// 16'hb5af, 16'hc071, 16'hcc7b, 16'hd994,
// 16'he770, 16'hf5cd, 16'h0462, 16'h12d9,
// 16'h20f8, 16'h2e62, 16'h3ae4, 16'h462d,
// 16'h5011, 16'h584e, 16'h5ecb, 16'h634e,
// 16'h65df, 16'h664f, 16'h64b9, 16'h6111,
// 16'h5b74, 16'h53fc, 16'h4ad1, 16'h4021,
// 16'h3425, 16'h271b, 16'h1944, 16'h0aec,
// 16'hfc5a, 16'heddc, 16'hdfbc, 16'hd243,
// 16'hc5b7, 16'hba59, 16'hb067, 16'ha80d,
// 16'ha182, 16'h9cda, 16'h9a3a, 16'h99a6,
// 16'h9b2a, 16'h9eb1, 16'ha43b, 16'hab97,
// 16'hb4b2, 16'hbf4c, 16'hcb3c, 16'hd838,
// 16'he608, 16'hf459, 16'h02ed, 16'h116a,
// 16'h1f94, 16'h2d16, 16'h39ae, 16'h451f,
// 16'h4f22, 16'h5793, 16'h5e35, 16'h62f9,
// 16'h65ad, 16'h6662, 16'h64f5, 16'h6188,
// 16'h5c18, 16'h54d1, 16'h4bcd, 16'h4144,
// 16'h3565, 16'h2871, 16'h1aaf, 16'h0c5e,
// 16'hfdd2, 16'hef49, 16'he122, 16'hd38f,
// 16'hc6ef, 16'hbb6a, 16'hb155, 16'ha8cf,
// 16'ha213, 16'h9d3b, 16'h9a65, 16'h999f,
// 16'h9ae8, 16'h9e44, 16'ha392, 16'haacb,
// 16'hb3b3, 16'hbe30, 16'hc9fa, 16'hd6e3,
// 16'he49e, 16'hf2e7, 16'h0177, 16'h0ffa,
// 16'h1e31, 16'h2bc3, 16'h387b, 16'h4407,
// 16'h4e35, 16'h56ce, 16'h5da1, 16'h6295,
// 16'h6580, 16'h6669, 16'h652f, 16'h61f9,
// 16'h5cb8, 16'h559f, 16'h4cc9, 16'h425e,
// 16'h36a5, 16'h29c8, 16'h1c15, 16'h0dd2,
// 16'hff45, 16'hf0bd, 16'he284, 16'hd4e4,
// 16'hc822, 16'hbc86, 16'hb242, 16'ha999,
// 16'ha2a6, 16'h9da4, 16'h9a93, 16'h999c,
// 16'h9ab0, 16'h9dd5, 16'ha2f7, 16'ha9fb,
// 16'hb2be, 16'hbd10, 16'hc8c3, 16'hd58a,
// 16'he33a, 16'hf173, 16'h2001, 16'h0e8a,
// 16'h1cca, 16'h2a72, 16'h3740, 16'h42ee,
// 16'h4d43, 16'h5604, 16'h5d0b, 16'h6228,
// 16'h6552, 16'h6663, 16'h656e, 16'h625c,
// 16'h5d59, 16'h5668, 16'h4dbd, 16'h437b,
// 16'h37de, 16'h2b1a, 16'h1d7f, 16'h0f41,
// 16'h20bc, 16'hf22e, 16'he3ea, 16'hd638,
// 16'hc95e, 16'hbd9d, 16'hb33b, 16'haa60,
// 16'ha346, 16'h9e0b, 16'h9acb, 16'h999c,
// 16'h9a7d, 16'h9d6d, 16'ha25e, 16'ha931,
// 16'hb1cd, 16'hbbf7, 16'hc788, 16'hd43a,
// 16'he1d1, 16'hf005, 16'hfe8a, 16'h0d18,
// 16'h1b63, 16'h291c, 16'h3606, 16'h41d0,
// 16'h4c4d, 16'h5537, 16'h5c6b, 16'h61bd,
// 16'h6518, 16'h6660, 16'h659e, 16'h62c2,
// 16'h5def, 16'h572f, 16'h4eae, 16'h4492,
// 16'h3915, 16'h2c6d, 16'h1ee3, 16'h10b1,
// 16'h0234, 16'hf39e, 16'he554, 16'hd78d,
// 16'hca9a, 16'hbebf, 16'hb431, 16'hab31,
// 16'ha3e6, 16'h9e7a, 16'h9b08, 16'h99a2,
// 16'h9a4e, 16'h9d0c, 16'ha1c7, 16'ha86f,
// 16'hb0dd, 16'hbae1, 16'hc653, 16'hd2e8,
// 16'he06e, 16'hee94, 16'hfd15, 16'h0ba5,
// 16'h19fa, 16'h27c6, 16'h34c6, 16'h40b2,
// 16'h4b50, 16'h5467, 16'h5bc7, 16'h614c,
// 16'h64d9, 16'h6659, 16'h65c6, 16'h6325,
// 16'h5e80, 16'h57f1, 16'h4f9b, 16'h45a6,
// 16'h3a49, 16'h2dbd, 16'h2045, 16'h1223,
// 16'h03a7, 16'hf513, 16'he6bc, 16'hd8e5,
// 16'hcbdc, 16'hbfde, 16'hb530, 16'hac02,
// 16'ha48d, 16'h9eee, 16'h9b4a, 16'h99ad,
// 16'h9a25, 16'h9cae, 16'ha137, 16'ha7b2,
// 16'hafef, 16'hb9d2, 16'hc51e, 16'hd19b,
// 16'hdf0c, 16'hed23, 16'hfba0, 16'h0a33,
// 16'h188e, 16'h266f, 16'h3383, 16'h3f8f,
// 16'h4a52, 16'h538f, 16'h5b21, 16'h60d5,
// 16'h6494, 16'h664c, 16'h65eb, 16'h6381,
// 16'h5f0d, 16'h58ae, 16'h5084, 16'h46b6,
// 16'h3b7a, 16'h2f0b, 16'h21a5, 16'h1394,
// 16'h051b, 16'hf686, 16'he829, 16'hda3c,
// 16'hcd22, 16'hc120, 16'hb632, 16'hacdc,
// 16'ha534, 16'h9f6b, 16'h9b8d, 16'h99c0,
// 16'h9a02, 16'h9c54, 16'ha0ae, 16'ha6f5,
// 16'haf0a, 16'hb8c4, 16'hc3ed, 16'hd050,
// 16'hddaa, 16'hebb5, 16'hfa2d, 16'h08bc,
// 16'h1726, 16'h2511, 16'h3240, 16'h3e69,
// 16'h494e, 16'h52b7, 16'h5a73, 16'h6058,
// 16'h644d, 16'h6635, 16'h6611, 16'h63d2,
// 16'h5f99, 16'h5963, 16'h516b, 16'h47c1,
// 16'h3caa, 16'h3054, 16'h2307, 16'h1520,
// 16'h0690, 16'hf7fc, 16'he992, 16'hdb9b,
// 16'hce65, 16'hc229, 16'hb738, 16'hadb5,
// 16'ha5e7, 16'h9fe6, 16'h9bda, 16'h99d7,
// 16'h99e2, 16'h9c01, 16'ha02a, 16'ha63c,
// 16'hae2b, 16'hb7b4, 16'hc2c5, 16'hcf04,
// 16'hdc4e, 16'hea44, 16'hf8ba, 16'h0746,
// 16'h15bb, 16'h23b4, 16'h30f9, 16'h3d3f,
// 16'h4848, 16'h51d7, 16'h59c3, 16'h5fd7,
// 16'h6420, 16'h661b, 16'h662c, 16'h6424,
// 16'h601a, 16'h5a1c, 16'h5247, 16'h48cc,
// 16'h3dd4, 16'h319c, 16'h2465, 16'h166d,
// 16'h0806, 16'hf96f, 16'heaff, 16'hdcfb,
// 16'hcfaa, 16'hc357, 16'hb83e, 16'hae98,
// 16'ha699, 16'ha06b, 16'h9c29, 16'h99f3,
// 16'h99c8, 16'h9bb7, 16'h9fa3, 16'ha590,
// 16'had47, 16'hb6b3, 16'hc198, 16'hcdbf,
// 16'hdaee, 16'he8db, 16'hf743, 16'h05d5,
// 16'h144a, 16'h2256, 16'h2fb0, 16'h3c12,
// 16'h473e, 16'h50f4, 16'h590d, 16'h5f51,
// 16'h63ac, 16'h65fe, 16'h6641, 16'h6470,
// 16'h6099, 16'h5ac9, 16'h5326, 16'h49cd,
// 16'h3f20, 16'h32de, 16'h25c5, 16'h17d6,
// 16'h097b, 16'hfae3, 16'hec6e, 16'hde5b,
// 16'hd0f4, 16'hc487, 16'hb948, 16'haf7e,
// 16'ha751, 16'ha0f3, 16'h9c81, 16'h9a12,
// 16'h99b6, 16'h9b6b, 16'h9f2a, 16'ha4e3,
// 16'hac6d, 16'hb5b0, 16'hc070, 16'hcc7c,
// 16'hd994, 16'he76f, 16'hf5cf, 16'h045f,
// 16'h12dd, 16'h20f4, 16'h2e66, 16'h3ae0,
// 16'h4631, 16'h500d, 16'h5853, 16'h5ec5,
// 16'h6354, 16'h65da, 16'h6652, 16'h64b9,
// 16'h610f, 16'h5b75, 16'h53fd, 16'h4acf,
// 16'h4024, 16'h3422, 16'h271d, 16'h1942,
// 16'h0aef, 16'hfc57, 16'heddf, 16'hdfba,
// 16'hd243, 16'hc5b8, 16'hba58, 16'hb067,
// 16'ha80f, 16'ha17f, 16'h9cdd, 16'h9a37,
// 16'h99a9, 16'h9b27, 16'h9eb4, 16'ha439,
// 16'hab98, 16'hb4b2, 16'hbf4b, 16'hcb3d,
// 16'hd838, 16'he608, 16'hf459, 16'h02ec,
// 16'h116b, 16'h1f93, 16'h2d18, 16'h39ab,
// 16'h4523, 16'h4f1e, 16'h5795, 16'h5e36,
// 16'h62f5, 16'h65b3, 16'h665d, 16'h64f8,
// 16'h6187, 16'h5c18, 16'h54d2, 16'h4bcb,
// 16'h4146, 16'h3563, 16'h2873, 16'h1aaf,
// 16'h0c5d, 16'hfdd1, 16'hef4c, 16'he11e,
// 16'hd394, 16'hc6e9, 16'hbb70, 16'hb150,
// 16'ha8d3, 16'ha20f, 16'h9d3f, 16'h9a62,
// 16'h99a1, 16'h9ae7, 16'h9e43, 16'ha395,
// 16'haac8, 16'hb3b6, 16'hbe2c, 16'hc9fe,
// 16'hd6e1, 16'he49f, 16'hf2e7, 16'h0174,
// 16'h0fff, 16'h1e2c, 16'h2bc7, 16'h3879,
// 16'h4406, 16'h4e38, 16'h56ca, 16'h5da5,
// 16'h6291, 16'h6584, 16'h6665, 16'h6533,
// 16'h61f5, 16'h5cbb, 16'h559e, 16'h4cc8,
// 16'h4261, 16'h36a1, 16'h29cb, 16'h1c13,
// 16'h0dd4, 16'hff44, 16'hf0bd, 16'he284,
// 16'hd4e3, 16'hc825, 16'hbc82, 16'hb246,
// 16'ha995, 16'ha2aa, 16'h9da1, 16'h9a96,
// 16'h9999, 16'h9ab2, 16'h9dd4, 16'ha2f7,
// 16'ha9fc, 16'hb2bc, 16'hbd14, 16'hc8be,
// 16'hd58e, 16'he337, 16'hf174, 16'h2002,
// 16'h0e89, 16'h1cca, 16'h2a73, 16'h373f,
// 16'h42f0, 16'h4d41, 16'h5605, 16'h5d0a,
// 16'h622a, 16'h6550, 16'h6666, 16'h6569,
// 16'h6261, 16'h5d55, 16'h566b, 16'h4dbb,
// 16'h437b, 16'h37df, 16'h2b1b, 16'h1d7c,
// 16'h0f44, 16'h20ba, 16'hf22e, 16'he3ed,
// 16'hd634, 16'hc95f, 16'hbda1, 16'hb335,
// 16'haa65, 16'ha344, 16'h9e09, 16'h9acf,
// 16'h999a, 16'h9a7d, 16'h9d6f, 16'ha25b,
// 16'ha934, 16'hb1ca, 16'hbbfa, 16'hc785,
// 16'hd43d, 16'he1cf, 16'hf006, 16'hfe89,
// 16'h0d1a, 16'h1b60, 16'h291f, 16'h3604,
// 16'h41d1, 16'h4c4d, 16'h5536, 16'h5c6c,
// 16'h61bd, 16'h6517, 16'h6662, 16'h659b,
// 16'h62c5, 16'h5ded, 16'h5730, 16'h4ead,
// 16'h4493, 16'h3915, 16'h2c6c, 16'h1ee4,
// 16'h10b1, 16'h0233, 16'hf39f, 16'he553,
// 16'hd78d, 16'hca9c, 16'hbebd, 16'hb431,
// 16'hab31, 16'ha3e6, 16'h9e7b, 16'h9b07,
// 16'h99a3, 16'h9a4d, 16'h9d0c, 16'ha1c8,
// 16'ha86f, 16'hb0db, 16'hbae5, 16'hc64e,
// 16'hd2ed, 16'he06b, 16'hee94, 16'hfd16,
// 16'h0ba4, 16'h19fb, 16'h27c5, 16'h34c7,
// 16'h40b0, 16'h4b52, 16'h5466, 16'h5bc7,
// 16'h614d, 16'h64d7, 16'h665a, 16'h65c6,
// 16'h6326, 16'h5e7e, 16'h57f3, 16'h4f99,
// 16'h45a8, 16'h3a48, 16'h2dbe, 16'h2043,
// 16'h1226, 16'h03a3, 16'hf517, 16'he6b9,
// 16'hd8e7, 16'hcbdb, 16'hbfde, 16'hb530,
// 16'hac02, 16'ha48e, 16'h9eed, 16'h9b4a,
// 16'h99ae, 16'h9a24, 16'h9caf, 16'ha138,
// 16'ha7af, 16'haff1, 16'hb9d1, 16'hc51f,
// 16'hd19b, 16'hdf0b, 16'hed24, 16'hfba0,
// 16'h0a32, 16'h188f, 16'h266e, 16'h3384,
// 16'h3f90, 16'h4a4f, 16'h5393, 16'h5b1d,
// 16'h60d8, 16'h6492, 16'h664d, 16'h65eb,
// 16'h6380, 16'h5f0e, 16'h58ae, 16'h5084,
// 16'h46b4, 16'h3b7d, 16'h2f09, 16'h21a7,
// 16'h1392, 16'h051c, 16'hf687, 16'he826,
// 16'hda41, 16'hcd1b, 16'hc107, 16'hb62e,
// 16'hacdc, 16'ha537, 16'h9f67, 16'h9b8f,
// 16'h99c0, 16'h9a20, 16'h9c58, 16'ha0aa,
// 16'ha6f8, 16'haf07, 16'hb8c6, 16'hc3ec,
// 16'hd050, 16'hddac, 16'hebb3, 16'hfa2d,
// 16'h08bc, 16'h1727, 16'h2510, 16'h3242,
// 16'h3e67, 16'h494f, 16'h52b6, 16'h5a75,
// 16'h6056, 16'h644f, 16'h6635, 16'h660e,
// 16'h63d6, 16'h5f96, 16'h5966, 16'h5169,
// 16'h47c1, 16'h3caa, 16'h3054, 16'h2307,
// 16'h1520, 16'h0691, 16'hf7fa, 16'he993,
// 16'hdb9b, 16'hce64, 16'hc22c, 16'hb734,
// 16'hadb8, 16'ha5e5, 16'h9fe8, 16'h9bd9,
// 16'h99d6, 16'h99e3, 16'h9c02, 16'ha027,
// 16'ha641, 16'hae24, 16'hb7bc, 16'hc2be,
// 16'hcf08, 16'hdc4c, 16'hea46, 16'hf8b9,
// 16'h0747, 16'h15b9, 16'h23b5, 16'h30f9,
// 16'h3d40, 16'h4846, 16'h51da, 16'h59bf,
// 16'h5fdb, 16'h63fc, 16'h661e, 16'h662a,
// 16'h6426, 16'h6019, 16'h5a1c, 16'h5246,
// 16'h48cd, 16'h3dd4, 16'h319d, 16'h2463,
// 16'h166f, 16'h0804, 16'hf971, 16'heafe,
// 16'hdcfb, 16'hcfa9, 16'hc35a, 16'hb83b,
// 16'hae9a, 16'ha698, 16'ha06b, 16'h9c2a,
// 16'h99f2, 16'h99c9, 16'h9bb6, 16'h9fa3,
// 16'ha592, 16'had44, 16'hb6b7, 16'hc193,
// 16'hcdc3, 16'hdaec, 16'he8dc, 16'hf743,
// 16'h05d4, 16'h144a, 16'h2257, 16'h2fb0,
// 16'h3c11, 16'h473f, 16'h50f3, 16'h590e,
// 16'h5f51, 16'h63ab, 16'h65ff, 16'h6640,
// 16'h6472, 16'h6098, 16'h5ac9, 16'h5325,
// 16'h49cf, 16'h3efe, 16'h32e1, 16'h25c1,
// 16'h17d9, 16'h0979, 16'hfae4, 16'hec70,
// 16'hde55, 16'hd0fc, 16'hc47f, 16'hb94e,
// 16'haf7b, 16'ha752, 16'ha0f3, 16'h9c80,
// 16'h9a13, 16'h99b5, 16'h9b6d, 16'h9f29,
// 16'ha4e2, 16'hac6d, 16'hb5b2, 16'hc06e,
// 16'hcc7e, 16'hd991, 16'he772, 16'hf5cc,
// 16'h0462, 16'h12da, 16'h20f7, 16'h2e63,
// 16'h3ae3, 16'h462d, 16'h5012, 16'h584e,
// 16'h5ec9, 16'h6351, 16'h65dd, 16'h6650,
// 16'h64b8, 16'h6112, 16'h5b72, 16'h53ff,
// 16'h4ace, 16'h4023, 16'h3425, 16'h271a,
// 16'h1945, 16'h0aeb, 16'hfc5b, 16'heddc,
// 16'hdfbc, 16'hd243, 16'hc5b6, 16'hba5b,
// 16'hb064, 16'ha810, 16'ha17f, 16'h9cdd,
// 16'h9a37, 16'h99a9, 16'h9b27, 16'h9eb4,
// 16'ha438, 16'hab9a, 16'hb4af, 16'hbf4f,
// 16'hcb3a, 16'hd839, 16'he607, 16'hf45a,
// 16'h02eb, 16'h116c, 16'h1f94, 16'h2d15,
// 16'h39af, 16'h451e, 16'h4f23, 16'h5792,
// 16'h5e37, 16'h62f6, 16'h65b1, 16'h665f,
// 16'h64f6, 16'h6189, 16'h5c16, 16'h54d3,
// 16'h4bcb, 16'h4146, 16'h3563, 16'h2873,
// 16'h1aae, 16'h0c5e, 16'hfdd2, 16'hef49,
// 16'he122, 16'hd38f, 16'hc6ee, 16'hbb6c,
// 16'hb153, 16'ha8d1, 16'ha212, 16'h9d3a,
// 16'h9a67, 16'h999c, 16'h9aec, 16'h9e40,
// 16'ha397, 16'haac6, 16'hb3b7, 16'hbe2c,
// 16'hc9fe, 16'hd6e0, 16'he4a0, 16'hf2e7,
// 16'h0174, 16'h0fff, 16'h1e2b, 16'h2bc8,
// 16'h3879, 16'h4406, 16'h4e37, 16'h56cc,
// 16'h5da3, 16'h6294, 16'h6581, 16'h6667,
// 16'h6531, 16'h61f8, 16'h5cb8, 16'h55a1,
// 16'h4cc5, 16'h4262, 16'h36a2, 16'h29c9,
// 16'h1c16, 16'h0dd1, 16'hff44, 16'hf0bf,
// 16'he282, 16'hd4e5, 16'hc823, 16'hbc84,
// 16'hb244, 16'ha997, 16'ha2a7, 16'h9da5,
// 16'h9a91, 16'h999f, 16'h9aad, 16'h9dd6,
// 16'ha2f8, 16'ha9f9, 16'hb2c0, 16'hbd10,
// 16'hc8c1, 16'hd58c, 16'he338, 16'hf175,
//  
//};
//assign depth = 44100; // same as numbers of row
///* end sine 1000 hz*/



/* shoot sound*/
 // stroe the value
logic [0:4079][15:0] ROM ={ // need to be 0 to 102 so first 2 bytes be on the left 
16'hFE3B, 16'hE468, 16'hE5E2, 16'h24F5,
 16'h5529, 16'h00BE, 16'h9E58, 16'hE894,
 16'h4B7D, 16'hF674, 16'hB69A, 16'hDB58,
 16'h0BB5, 16'h603E, 16'h17CE, 16'hBD27,
 16'hD2E3, 16'h1A14, 16'h37F5, 16'hE502,
 16'hCB06, 16'h00F3, 16'h5013, 16'h06EA,
 16'hAE18, 16'hDDE6, 16'hFC1C, 16'h4EE2,
 16'h251F, 16'hC7E2, 16'hCE1C, 16'h06E7,
 16'h4215, 16'hF4F0, 16'hC40A, 16'hF8FD,
 16'h4CFA, 16'h070F, 16'hBFE9, 16'hEA20,
 16'h0ED6, 16'h2C34, 16'hE8C1, 16'hB54A,
 16'hF9AB, 16'h4760, 16'h0496, 16'hCA73,
 16'hE885, 16'h5782, 16'h6A77, 16'hDB8F,
 16'hA96D, 16'hD495, 16'h226A, 16'hF296,
 16'hA16B, 16'hD094, 16'h156D, 16'h5090,
 16'h3774, 16'h4589, 16'h3E7A, 16'hF083,
 16'hDE7E, 16'h8C82, 16'h8000, 16'hCF83,
 16'h257B, 16'hEF89, 16'hF771, 16'h6E96,
 16'h7D63, 16'h7FA4, 16'hF455, 16'h80B2,
 16'h8000, 16'h80C0, 16'h8000, 16'h80C3,
 16'hD73F, 16'h6CBC, 16'h7D4C, 16'h7FAA,
 16'h7D65, 16'h7F86, 16'h3C92, 16'h8053,
 16'h8000, 16'h800D, 16'h931B, 16'h29B8,
 16'h2178, 16'h0757, 16'h7FDC, 16'h7CEF,
 16'h7FFF, 16'h3284, 16'hA6AF, 16'h8001,
 16'h8210, 16'h8CC2, 16'h826B, 16'hB96B,
 16'h28BB, 16'h7C23, 16'h7FFF, 16'h7BEA,
 16'h7FFF, 16'h7BBB, 16'hBE59, 16'h8000,
 16'h837A, 16'hA578, 16'hBE95, 16'hA85F,
 16'h03AD, 16'h4E48, 16'h7FFF, 16'h7A35,
 16'h7FFF, 16'h1228, 16'hB5DE, 16'h881D,
 16'h83E6, 16'h8000, 16'h8CE5, 16'h0420,
 16'h4CD7, 16'h4C35, 16'h6FBC, 16'h7A57,
 16'h7FFF, 16'h4C87, 16'h835B, 16'h8000,
 16'h8317, 16'h8B0E, 16'h92CD, 16'h9C59,
 16'h0180, 16'h7CA6, 16'h7FFC, 16'h7CEA,
 16'h7FFC, 16'h7A1A, 16'h11D5, 16'h8000,
 16'h81C2, 16'h8000, 16'hCDC0, 16'hC239,
 16'hCBD3, 16'h291D, 16'h7FFE, 16'h7CF3,
 16'h7FFE, 16'h66C5, 16'h0C51, 16'hB29B,
 16'h8276, 16'h8003, 16'h8A88, 16'hE777,
 16'hCF83, 16'hF88B, 16'h535F, 16'h7BBF,
 16'h7FFE, 16'h7C14, 16'h13B7, 16'hC185,
 16'h8837, 16'h8000, 16'h809E, 16'h8000,
 16'h06F5, 16'h2562, 16'h1E48, 16'h5B0D,
 16'h7D9E, 16'h7FB4, 16'h7CFD, 16'hD34F,
 16'h8000, 16'h82D7, 16'h8000, 16'h8345,
 16'h8000, 16'hD496, 16'h524C, 16'h63CB,
 16'h6125, 16'h7FFF, 16'h7B1A, 16'h7FFE,
 16'hEE28, 16'h83C8, 16'h8001, 16'h8393,
 16'hC78F, 16'hC149, 16'hABE5, 16'hFFE8,
 16'h4E50, 16'h7FFF, 16'h7CD0, 16'h7FE8,
 16'h5C63, 16'hF74E, 16'hB504, 16'h80AA,
 16'h8000, 16'h8007, 16'hF049, 16'h0369,
 16'hE7E1, 16'h36DA, 16'h7FFF, 16'h7D62,
 16'h7FFF, 16'h5B0D, 16'h0A0D, 16'hC6E5,
 16'h821D, 16'h8000, 16'h81F9, 16'hE42C,
 16'hE1A1, 16'hDFA0, 16'h3213, 16'h7D44,
 16'h7F5B, 16'h7E0F, 16'h7E81, 16'h3EF4,
 16'hF593, 16'h81E8, 16'h8001, 16'h82DE,
 16'hA8AB, 16'hFFC7, 16'hEFCE, 16'hFD93,
 16'h5917, 16'h7FFF, 16'h7990, 16'h7FFF,
 16'h6545, 16'hE7CA, 16'hAB35, 16'h85BD,
 16'h8000, 16'h8576, 16'h8AC3, 16'h05F8,
 16'h4A57, 16'h2852, 16'h3D0B, 16'h7FFF,
 16'h7AD5, 16'h7FFF, 16'h43AA, 16'h93EA,
 16'h8000, 16'h811B, 16'h8002, 16'h8062,
 16'hA7EE, 16'h19CA, 16'h4C75, 16'h3E57,
 16'h50D3, 16'h7E0C, 16'h7F0B, 16'h7DE9,
 16'h141A, 16'hC8EB, 16'h9407, 16'h8000,
 16'h80D5, 16'h8001, 16'hEF92, 16'h0B93,
 16'hF746, 16'h33E3, 16'h7EF5, 16'h7E30,
 16'h7EAE, 16'h6B70, 16'h5177, 16'hFA9E,
 16'h8000, 16'h80BA, 16'h8000, 16'hA1BA,
 16'hD350, 16'hD19F, 16'hF978, 16'h4F6C,
 16'h7DB4, 16'h7F28, 16'h7DFF, 16'h7ED8,
 16'h7F52, 16'h0283, 16'h80A7, 16'h8001,
 16'h80F7, 16'h9BE5, 16'h9F3A, 16'h9FAA,
 16'hF36D, 16'h3683, 16'h7F87, 16'h7D75,
 16'h7988, 16'h7D82, 16'h7F6D, 16'h60AA,
 16'hA239, 16'h8001, 16'h80ED, 16'h8000,
 16'hB78B, 16'hABAC, 16'hB91A, 16'h0022,
 16'h559F, 16'h7FA2, 16'h721D, 16'h7F23,
 16'h7D9F, 16'h7F9C, 16'h602A, 16'hA50F,
 16'h8003, 16'h8278, 16'h8000, 16'h8ECE,
 16'h9C10, 16'hE40D, 16'h26DB, 16'h6B38,
 16'h5CBB, 16'h674C, 16'h7AB3, 16'h7FFE,
 16'h7BC3, 16'h0F2E, 16'hA2E7, 16'h82FF,
 16'h8000, 16'h82BE, 16'h8000, 16'h8E6B,
 16'hDDC3, 16'h410C, 16'h3E27, 16'h2EA5,
 16'h7090, 16'h7FFF, 16'h7CFA, 16'h7FD3,
 16'h4D5E, 16'hB274, 16'h8004, 16'h8023,
 16'h8003, 16'h8000, 16'h8034, 16'hC5B7,
 16'h1459, 16'h679C, 16'h3F6A, 16'h3E96,
 16'h7766, 16'h7EA1, 16'h7F56, 16'h6AB3,
 16'h0C42, 16'hA6CC, 16'h8025, 16'h8000,
 16'h8005, 16'h8009, 16'h96EB, 16'hF61F,
 16'h4EDA, 16'h272B, 16'h22D2, 16'h5F2E,
 16'h7ED5, 16'h7E25, 16'h7EE4, 16'h5110,
 16'h07FE, 16'hBEF4, 16'h891A, 16'h8000,
 16'h8037, 16'h8000, 16'hD74C, 16'hF7AE,
 16'hF254, 16'h18AD, 16'h344F, 16'h7BB8,
 16'h7F3D, 16'h7DD2, 16'h641C, 16'h6DF9,
 16'h5AEF, 16'hD62C, 16'h8000, 16'h8068,
 16'h8000, 16'h80A6, 16'h943E, 16'hB6DE,
 16'h0106, 16'h4C14, 16'h46D3, 16'h3145,
 16'h6CA7, 16'h7F69, 16'h7D8A, 16'h677F,
 16'h4E7C, 16'h0987, 16'hC978, 16'h8187,
 16'h8002, 16'h8183, 16'h8002, 16'hDF7F,
 16'hE682, 16'hF17E, 16'h2F80, 16'h6283,
 16'h4979, 16'h588E, 16'h7D69, 16'h7FA1,
 16'h7D53, 16'h49BA, 16'hEE38, 16'hACD7,
 16'h8819, 16'h81F8, 16'h8000, 16'h8218,
 16'hD8DB, 16'hE62E, 16'hF0CE, 16'h2832,
 16'h53D2, 16'h7626, 16'h65E5, 16'h5A0B,
 16'h7D0B, 16'h7FDA, 16'h5F46, 16'h1696,
 16'hBD91, 16'h9745, 16'h8000, 16'h80E7,
 16'h8000, 16'hA783, 16'hE4B0, 16'hF01D,
 16'h0C14, 16'h44BD, 16'h5870, 16'h4467,
 16'h5BBC, 16'h7D25, 16'h7FF6, 16'h66F4,
 16'h351D, 16'h07D8, 16'hD12D, 16'h8FD3,
 16'h8127, 16'h8000, 16'h810D, 16'hBE06,
 16'hCEE2, 16'hEB39, 16'h19AB, 16'h4473,
 16'h706F, 16'h52AE, 16'h4F35, 16'h67E7,
 16'h7EFF, 16'h7E19, 16'h50D3, 16'h0F3C,
 16'hC6B8, 16'hA450, 16'h8000, 16'h8050,
 16'h8000, 16'h963F, 16'hE5D1, 16'hEA1C,
 16'h06FB, 16'h29EA, 16'h4833, 16'h77AE,
 16'h5D74, 16'h5368, 16'h69BC, 16'h7D20,
 16'h7FFF, 16'h41DE, 16'hF03E, 16'hA3A9,
 16'h866E, 16'h8001, 16'h8193, 16'h8000,
 16'h9BA6, 16'hFC59, 16'h00A3, 16'h0964,
 16'h2D90, 16'h3C81, 16'h606B, 16'h71AD,
 16'h5D37, 16'h54E7, 16'h69F9, 16'h7D29,
 16'h5DB5, 16'h0E6D, 16'hB671, 16'h81B0,
 16'h8030, 16'h8000, 16'h8001, 16'h8025,
 16'hC1C3, 16'h1A53, 16'h2F99, 16'h2178,
 16'h2B7A, 16'h2B92, 16'h5464, 16'h7AA4,
 16'h5C55, 16'h52B0, 16'h604E, 16'h73B3,
 16'h4A4C, 16'hFAB4, 16'hAE4D, 16'h89B2,
 16'h8150, 16'h80AD, 16'h8001, 16'h82A9,
 16'hCA58, 16'h19A8, 16'h2658, 16'h1FA8,
 16'h3058, 16'h4AA7, 16'h585A, 16'h43A6,
 16'h415A, 16'h5DA6, 16'h7759, 16'h6BA7,
 16'h3A5A, 16'h0FA3, 16'hE862, 16'hB499,
 16'h8000, 16'h808C, 16'h8001, 16'h8F7D,
 16'hBE8D, 16'hCE6B, 16'h049C, 16'h265C,
 16'h48AB, 16'h5750, 16'h2CB5, 16'h2047,
 16'h3DBC, 16'h7040, 16'h63C3, 16'h4D3C,
 16'h47C4, 16'h4E3F, 16'h4BBC, 16'hEC49,
 16'h93B1, 16'h8057, 16'h8000, 16'h8068,
 16'h8001, 16'h9280, 16'hD875, 16'h2397,
 16'h2D5D, 16'h22AC, 16'h274D, 16'h3ABA,
 16'h5740, 16'h36C4, 16'h2A3B, 16'h49C3,
 16'h5241, 16'h70B9, 16'h524F, 16'h2BA7,
 16'h1866, 16'hF189, 16'hC28C, 16'h805D,
 16'h8000, 16'h802B, 16'h8001, 16'h8EF2,
 16'hB52B, 16'hF2B8, 16'h1763, 16'h4784,
 16'h5595, 16'h3153, 16'h1DC3, 16'h2F29,
 16'h48E8, 16'h3F0B, 16'h3100, 16'h41F8,
 16'h5A0C, 16'h4EF3, 16'h290C, 16'h05F8,
 16'hD801, 16'hB509, 16'h82EA, 16'h8000,
 16'h80C9, 16'h8000, 16'hB6A0, 16'hCC77,
 16'hEB72, 16'h17A4, 16'h3446, 16'h52D0,
 16'h451B, 16'h25FA, 16'h28F1, 16'h3B23,
 16'h41CB, 16'h3545, 16'h38AE, 16'h4C5D,
 16'h599A, 16'h2D6E, 16'h148A, 16'h037D,
 16'hDA7E, 16'hBC85, 16'h8000, 16'h8086,
 16'h8000, 16'h8282, 16'hBF81, 16'hD77C,
 16'hEB87, 16'h1F76, 16'h448E, 16'h456D,
 16'h3398, 16'h2764, 16'h30A0, 16'h415B,
 16'h2CA9, 16'h1F53, 16'h36B2, 16'h3E49,
 16'h55BD, 16'h493A, 16'h1FD0, 16'h1827,
 16'h0BE0, 16'hE61A, 16'hA1EC, 16'h800D,
 16'h8000, 16'h81FB, 16'h860E, 16'h91E9,
 16'hC721, 16'hF2D5, 16'h2534, 16'h4BC4,
 16'h3744, 16'h29B4, 16'h3754, 16'h43A4,
 16'h2664, 16'h0F96, 16'h176D, 16'h3390,
 16'h4C74, 16'h4089, 16'h2E7A, 16'h3283,
 16'h397E, 16'h1C82, 16'h037E, 16'hDF83,
 16'hBB7C, 16'hA384, 16'h807C, 16'h8001,
 16'h807C, 16'h9684, 16'hCE7B, 16'hE784,
 16'hFD7E, 16'h1A80, 16'h3983, 16'h4979,
 16'h308B, 16'h2771, 16'h2793, 16'h3469,
 16'h299B, 16'h0D61, 16'h19A4, 16'h3357,
 16'h49AD, 16'h334F, 16'h27B4, 16'h274A,
 16'h2AB8, 16'h2946, 16'h00BB, 16'hD346,
 16'hACB7, 16'h9D4E, 16'h8FAB, 16'h8005,
 16'h829D, 16'h956B, 16'hBA8C, 16'hF67F,
 16'h0972, 16'h149F, 16'h2C50, 16'h2FC2,
 16'h422C, 16'h38E5, 16'h2409, 16'h1B09,
 16'h1BE6, 16'h292B, 16'h11C4, 16'h074C,
 16'h20A5, 16'h3869, 16'h3E8C, 16'h2B7D,
 16'h1B7C, 16'h2289, 16'h2774, 16'h0E8D,
 16'hEB76, 16'hD484, 16'hBB84, 16'h9072,
 16'h8003, 16'h875D, 16'h9CAE, 16'hB046,
 16'hB5C7, 16'hD52B, 16'hFFE4, 16'h2A0D,
 16'h3703, 16'h29ED, 16'h3222, 16'h39D1,
 16'h313A, 16'h1FBD, 16'h124A, 16'h16B1,
 16'h2053, 16'h10AB, 16'h0555, 16'h14AC,
 16'h2752, 16'h3BB1, 16'h294B, 16'h19BC,
 16'h1E3B, 16'h1ECE, 16'h1C28, 16'h01E3,
 16'hED13, 16'hDFF6, 16'hC401, 16'h9708,
 16'h84F1, 16'h8D15, 16'h96E5, 16'hB220,
 16'hC6DD, 16'hD024, 16'hE9DE, 16'h111E,
 16'h27E6, 16'h3B15, 16'h3EF2, 16'h2D06,
 16'h2A03, 16'h27F2, 16'h2D1A, 16'h20DB,
 16'h0A2E, 16'h0ACA, 16'h133D, 16'h0EBE,
 16'h0447, 16'h0CB4, 16'h1F4E, 16'h2FB2,
 16'h2D4D, 16'h1EB7, 16'h1942, 16'h14C6,
 16'h1330, 16'h15DD, 16'hFF15, 16'hECFA,
 16'hDAF4, 16'hB420, 16'hABCB, 16'hA14B,
 16'h8E9F, 16'h9776, 16'hA776, 16'hC59D,
 16'hD150, 16'hDFC2, 16'hFD2D, 16'h14E2,
 16'h3313, 16'h37F5, 16'h3105, 16'h2CFF,
 16'h2CFF, 16'h3101, 16'h2502, 16'h0FF8,
 16'h0F12, 16'h14E0, 16'h1530, 16'h09BF,
 16'hFD53, 16'h009B, 16'h0E77, 16'h1474,
 16'h18A3, 16'h1C47, 16'h21CE, 16'h281F,
 16'h13F1, 16'h0B00, 16'h070E, 16'h06E5,
 16'h0727, 16'hF5CF, 16'hE939, 16'hDBC1,
 16'hC942, 16'hADBE, 16'h9940, 16'h9EC5,
 16'hAC33, 16'hB5D7, 16'hBC1E, 16'hC9EE,
 16'hDB06, 16'hF606, 16'h11ED, 16'h1B21,
 16'h25D0, 16'h2D3F, 16'h35B3, 16'h375A,
 16'h279A, 16'h2170, 16'h1E87, 16'h1E81,
 16'h1B79, 16'h0D8B, 16'h0A72, 16'h0E8F,
 16'h0E72, 16'h038C, 16'hFF77, 16'h0184,
 16'h0A82, 16'h0F77, 16'h0892, 16'h0E64,
 16'h17A5, 16'h2252, 16'h1FB8, 16'h133E,
 16'h0ACD, 16'h0527, 16'h06E4, 16'h0113,
 16'hF2F5, 16'hF004, 16'hF502, 16'hEEFA,
 16'hD907, 16'hC2F9, 16'hB205, 16'hACFF,
 16'hB4FC, 16'hB40A, 16'hB9EF, 16'hC21A,
 16'hD3DB, 16'hE931, 16'hE7C2, 16'hF14C,
 16'h06A7, 16'h1C65, 16'h288F, 16'h2B7E,
 16'h2C75, 16'h2F98, 16'h305B, 16'h26B1,
 16'h1F45, 16'h18C3, 16'h1737, 16'h18CF,
 16'h0B2B, 16'h0ADA, 16'h0D23, 16'h0BDE,
 16'h0B23, 16'h01DA, 16'h032A, 16'h00D2,
 16'h0833, 16'h04C8, 16'hFF3D, 16'hFFBD,
 16'h0649, 16'h0BB1, 16'h0D55, 16'h0FA6,
 16'h115F, 16'h169B, 16'h106B, 16'h088F,
 16'h0175, 16'h008A, 16'hFD76, 16'h008A,
 16'hF277, 16'hEF86, 16'hF07F, 16'hF77B,
 16'hF68C, 16'hD66C, 16'hAD9C, 16'h8C5C,
 16'h8000, 16'h8646, 16'hB3C9, 16'hE025,
 16'h0AEF, 16'h1FFD, 16'h4817, 16'h7ED4,
 16'h7E42, 16'h2DA8, 16'hD16E, 16'hB97C,
 16'hB69A, 16'hE751, 16'h5BC2, 16'h4E2D,
 16'hD2E1, 16'hC614, 16'hC5F5, 16'hEF04,
 16'h6C00, 16'h49FF, 16'hD000, 16'hC404,
 16'hC7F4, 16'hF718, 16'h6ED8, 16'h4E3B,
 16'hCFB0, 16'hC267, 16'hC381, 16'hF498,
 16'h724D, 16'h4ACE, 16'hCE18, 16'hC002,
 16'hBFE6, 16'hF02F, 16'h70BE, 16'h4F52,
 16'hCDA1, 16'hBF69, 16'hBB91, 16'hEC72,
 16'h728E, 16'h526E, 16'hCC98, 16'hBA5E,
 16'hB7B1, 16'hE73D, 16'h73D7, 16'h5812,
 16'hD106, 16'hBAE1, 16'hBA39, 16'hE1AD,
 16'h686C, 16'h5F7B, 16'hD29D, 16'hB34E,
 16'hBAC4, 16'hD62D, 16'h5DDF, 16'h6B18,
 16'hE1ED, 16'hB413, 16'hB9E8, 16'hD022,
 16'h4CD0, 16'h7941, 16'hF5AB, 16'hB26D,
 16'hB676, 16'hC7AB, 16'h3632, 16'h7EF3,
 16'h09E7, 16'hB33E, 16'hB89E, 16'hBE86,
 16'h2657, 16'h7ECA, 16'h2317, 16'hB706,
 16'hB4E1, 16'hB932, 16'h0DC1, 16'h7F45,
 16'h3DBC, 16'hBB3D, 16'hB2D0, 16'hB81D,
 16'hF1FA, 16'h7FEB, 16'h5435, 16'hCBA6,
 16'hB285, 16'hB64B, 16'hDFE9, 16'h66E1,
 16'h7355, 16'hDF75, 16'hABC2, 16'hB508,
 16'hCE2B, 16'h46A5, 16'h7FFF, 16'h0353,
 16'hAFCE, 16'hB717, 16'hBFFE, 16'h20F4,
 16'h7FFF, 16'h2EF0, 16'hB608, 16'hB508,
 16'hB8E1, 16'hF73D, 16'h7FFF, 16'h548F,
 16'hC140, 16'hADF5, 16'hB2D4, 16'hE165,
 16'h6D5F, 16'h74DE, 16'hE0E6, 16'hAE55,
 16'hBA72, 16'hCBC3, 16'h3D0D, 16'h7FFF,
 16'h13BD, 16'hAF62, 16'hB284, 16'hB891,
 16'h0C60, 16'h7FA9, 16'h4753, 16'hBAAB,
 16'hAE5C, 16'hB298, 16'hE378, 16'h7374,
 16'h71A4, 16'hDB41, 16'hAADC, 16'hB305,
 16'hC51A, 16'h3DC8, 16'h7E55, 16'h1791,
 16'hAD87, 16'hB562, 16'hB9B3, 16'h003A,
 16'h7ED8, 16'h531A, 16'hC3F0, 16'hAB09,
 16'hB1FB, 16'hDB03, 16'h5DFE, 16'h7F02,
 16'hF3FE, 16'hAA03, 16'hB5FA, 16'hBC0A,
 16'h23F1, 16'h7E13, 16'h3AEC, 16'hB313,
 16'hACEF, 16'hB50E, 16'hE5F4, 16'h780B,
 16'h75F8, 16'hDD03, 16'hA902, 16'hB5F8,
 16'hC010, 16'h2FE9, 16'h7E1E, 16'h2DDA,
 16'hAF2D, 16'hACCD, 16'hB63A, 16'hEFC0,
 16'h7F44, 16'h6AB8, 16'hD14A, 16'hA6B7,
 16'hB648, 16'hC6B9, 16'h3144, 16'h7EC0,
 16'h273B, 16'hAECB, 16'hAF2F, 16'hB9D7,
 16'hEE24, 16'h7BE1, 16'h7518, 16'hD7EF,
 16'hAE0A, 16'hB1FF, 16'hC6F8, 16'h3010,
 16'h7DE7, 16'h3422, 16'hB1D7, 16'hAD2F,
 16'hB5CA, 16'hE43D, 16'h6ABC, 16'h7E4B,
 16'hE9AF, 16'hA856, 16'hB5A5, 16'hC060,
 16'h179C, 16'h7E68, 16'h4E94, 16'hBE6F,
 16'hA68F, 16'hB273, 16'hD78C, 16'h4975,
 16'h7E89, 16'h0B79, 16'hA786, 16'hAF7B,
 16'hB685, 16'hF77A, 16'h7E87, 16'h7079,
 16'hD087, 16'hA87B, 16'hB381, 16'hC484,
 16'h2177, 16'h7F8E, 16'h3D6D, 16'hB398,
 16'hAC63, 16'hB2A3, 16'hDC57, 16'h56AD,
 16'h7E50, 16'h07B4, 16'hA748, 16'hB4BC,
 16'hB83F, 16'hF7C4, 16'h7E3D, 16'h71C0,
 16'hD745, 16'hA8B3, 16'hB555, 16'hC5A3,
 16'h1B67, 16'h7F8D, 16'h4E81, 16'hBB6E,
 16'hAAA5, 16'hB447, 16'hD4CF, 16'h3D1A,
 16'h7EFD, 16'h24EC, 16'hAE2A, 16'hAEC2,
 16'hBB51, 16'hE49D, 16'h5D72, 16'h7E82,
 16'hFC89, 16'hA86D, 16'hB09A, 16'hBB63,
 16'hFA9D, 16'h7D67, 16'h7391, 16'hDE79,
 16'hA57C, 16'hB192, 16'hC65E, 16'h0FB3,
 16'h7E39, 16'h5CDC, 16'hC210, 16'hA905,
 16'hB5E6, 16'hCA2C, 16'h23C4, 16'h7E4B,
 16'h47A8, 16'hB663, 16'hAA95, 16'hB46F,
 16'hD391, 16'h376C, 16'h7E9A, 16'h305E,
 16'hB1AD, 16'hAD44, 16'hB8CE, 16'hDE1E,
 16'h48F8, 16'h7DF2, 16'h1C24, 16'hAEC4,
 16'hAE55, 16'hBB92, 16'hE486, 16'h5764,
 16'h7FAE, 16'h0944, 16'hACC8, 16'hB02F,
 16'hBDD6, 16'hEF27, 16'h5FDA, 16'h7E2A,
 16'hFDCE, 16'hAB3D, 16'hB2B3, 16'hC060,
 16'hF08C, 16'h648A, 16'h7E5E, 16'hF8BB,
 16'hA72A, 16'hAEF1, 16'hBEF6, 16'hF322,
 16'h6AC7, 16'h7F4E, 16'hF79F, 16'hAE72,
 16'hAF81, 16'hBF88, 16'hF671, 16'h6693,
 16'h7E6D, 16'hF590, 16'hAA77, 16'hB17E,
 16'hC390, 16'hF35F, 16'h64B6, 16'h7E32,
 16'hFFE7, 16'hAE01, 16'hAE17, 16'hC2D1,
 16'hEF47, 16'h5AA0, 16'h7E79, 16'h0671,
 16'hAFA2, 16'hB34E, 16'hBFBF, 16'hEB38,
 16'h4CCF, 16'h7E2C, 16'h19D5, 16'hB12D,
 16'hAFCF, 16'hBC39, 16'hE1BB, 16'h3F52,
 16'h7E9E, 16'h2975, 16'hB178, 16'hB19A,
 16'hBA53, 16'hDAC0, 16'h2D2D, 16'h7DE6,
 16'h4308, 16'hB907, 16'hA5EE, 16'hAE1B,
 16'hCBDC, 16'h152C, 16'h7DCE, 16'h5036,
 16'hBFCA, 16'hA232, 16'hB1D4, 16'hCE24,
 16'h07E6, 16'h7F0F, 16'h68FC, 16'hCEF8,
 16'hA815, 16'hB1DE, 16'hC730, 16'hF6C2,
 16'h684B, 16'h7DA9, 16'hF062, 16'hAA94,
 16'hAE75, 16'hC283, 16'hE984, 16'h4876,
 16'h7F8E, 16'h1E6F, 16'hAF94, 16'hAD6A,
 16'hBC96, 16'hDA6B, 16'h2A94, 16'h7E6E,
 16'h4790, 16'hBE71, 16'hAD8E, 16'hB672,
 16'hD28F, 16'h0C70, 16'h7F90, 16'h7170,
 16'hDA90, 16'hAF6F, 16'hB193, 16'hCA6B,
 16'hF597, 16'h5367, 16'h7F9A, 16'h1166,
 16'hAF9A, 16'hAE66, 16'hBE9A, 16'hE467,
 16'h2697, 16'h7E6D, 16'h498C, 16'hBE7D,
 16'hAF79, 16'hB792, 16'hD462, 16'h06AB,
 16'h7347, 16'h7CC8, 16'hE927, 16'hABEA,
 16'hB705, 16'hC60C, 16'hEEE4, 16'h3C2A,
 16'h7DC9, 16'h3142, 16'hB5B6, 16'hAF4F,
 16'hB6AF, 16'hDA50, 16'h11B4, 16'h7B44,
 16'h72C8, 16'hDB26, 16'hAEF2, 16'hB5F1,
 16'hCC30, 16'hF0AD, 16'h3E77, 16'h7E63,
 16'h27C4, 16'hB516, 16'hB010, 16'hBDCA,
 16'hDD5B, 16'h0E81, 16'h7AA1, 16'h7141,
 16'hE0D7, 16'hB118, 16'hB3F2, 16'hC80B,
 16'hEAF1, 16'h361A, 16'h7FD3, 16'h3748,
 16'hB995, 16'hAE96, 16'hB638, 16'hD5FE,
 16'h05C8, 16'h6776, 16'h7F48, 16'hF2FE,
 16'hB1BA, 16'hB38E, 16'hBF2D, 16'hEA13,
 16'h21B2, 16'h7FFD, 16'h5448, 16'hC3E3,
 16'hADFA, 16'hB620, 16'hD1D0, 16'hF836,
 16'h45CD, 16'h7FFF, 16'h1DF3, 16'hB7EB,
 16'hB13F, 16'hBB8E, 16'hDDAD, 16'h0C13,
 16'h7133, 16'h7B81, 16'hEBCE, 16'hAFE2,
 16'hB26F, 16'hC241, 16'hE50C, 16'h1DA9,
 16'h7F9E, 16'h5620, 16'hC81D, 16'hAFAD,
 16'hB381, 16'hCE58, 16'hF3C7, 16'h3022,
 16'h7FFF, 16'h3709, 16'hBBF7, 16'hAC12,
 16'hB6DE, 16'hD539, 16'hFCAA, 16'h4976,
 16'h7FFF, 16'h16C3, 16'hB310, 16'hAE20,
 16'hBDAD, 16'hDE87, 16'h0746, 16'h60ED,
 16'h7EDF, 16'hFA55, 16'hB277, 16'hB4BD,
 16'hC012, 16'hE21B, 16'h0EB9, 16'h7272,
 16'h6E66, 16'hE6C0, 16'hAE1C, 16'hB104,
 16'hC5DF, 16'hE83D, 16'h10A9, 16'h7F6F,
 16'h667B, 16'hD499, 16'hB054, 16'hB5BD,
 16'hC835, 16'hE7D7, 16'h1A20, 16'h7FE6,
 16'h5C16, 16'hD4EC, 16'hB114, 16'hB6EC,
 16'hCD16, 16'hEAE6, 16'h1D1F, 16'h7FDA,
 16'h5E30, 16'hCEC5, 16'hB347, 16'hB7AB,
 16'hC864, 16'hEB8D, 16'h1882, 16'h7F6E,
 16'h60A3, 16'hD54C, 16'hB1C4, 16'hB72D,
 16'hC9E1, 16'hEA12, 16'h15FA, 16'h7FFB,
 16'h630F, 16'hD8E9, 16'hB21E, 16'hB5DB,
 16'hC92B, 16'hE9D0, 16'h1235, 16'h74C6,
 16'h6D3E, 16'hE9BE, 16'hB147, 16'hB1B3,
 16'hC954, 16'hE6A2, 16'h0A6A, 16'h6689,
 16'h7986, 16'hFD69, 16'hB4A9, 16'hB543,
 16'hBFD4, 16'hE513, 16'h0008, 16'h4FDB,
 16'h7E43, 16'h129D, 16'hB685, 16'hB359,
 16'hBDC8, 16'hD918, 16'hF907, 16'h3DDB,
 16'h7FFC, 16'h2EA2, 16'hBE78, 16'hAC72,
 16'hBA9F, 16'hD556, 16'hF3B0, 16'h224E,
 16'h7FAE, 16'h515B, 16'hC797, 16'hB47D,
 16'hB56A, 16'hCCB3, 16'hEE2B, 16'h10FB,
 16'h72DB, 16'h6F53, 16'hEB7E, 16'hB6B1,
 16'hB61F, 16'hC111, 16'hE7BF, 16'h0071,
 16'h4861, 16'h7FCA, 16'h1B0E, 16'hBA16,
 16'hB1CC, 16'hBA4C, 16'hE0A1, 16'hF46D,
 16'h288B, 16'h7FFF, 16'h4D8E, 16'hCB67,
 16'hB0AA, 16'hB63F, 16'hCCDC, 16'hF105,
 16'h0D1F, 16'h64BA, 16'h7B6F, 16'h0067,
 16'hB5C3, 16'hB313, 16'hBF16, 16'hE5C3,
 16'hFA63, 16'h3379, 16'h7FA6, 16'h413F,
 16'hC3DA, 16'hAE11, 16'hB9FE, 16'hD6F7,
 16'hF010, 16'h0DF0, 16'h690B, 16'h77FC,
 16'hFAF9, 16'hB915, 16'hB7DB, 16'hC237,
 16'hE6B4, 16'hF564, 16'h3082, 16'h7D98,
 16'h434F, 16'hC6C9, 16'hB321, 16'hB9F4,
 16'hD2F7, 16'hF01C, 16'h06D4, 16'h583B,
 16'h7DB8, 16'h1652, 16'hB5A6, 16'hB35F,
 16'hBB9F, 16'hDB62, 16'hF29E, 16'h1E61,
 16'h7CA1, 16'h645B, 16'hE2AB, 16'hB54D,
 16'hB9BC, 16'hC73A, 16'hE6D1, 16'hFA24,
 16'h31E6, 16'h7F11, 16'h41F7, 16'hC402,
 16'hB405, 16'hBBF4, 16'hD013, 16'hF0E6,
 16'h0720, 16'h4EDB, 16'h7E2A, 16'h23D2,
 16'hBD31, 16'hB1CB, 16'hBA38, 16'hD7C7,
 16'hF73A, 16'h0EC6, 16'h6138, 16'h7DC9,
 16'h0936, 16'hB8CD, 16'hB630, 16'hBED3,
 16'hDE29, 16'hF6DC, 16'h191F, 16'h6EE6,
 16'h6F16, 16'hEFEE, 16'hB50E, 16'hB9F6,
 16'hC406, 16'hE700, 16'hF6FA, 16'h1B0B,
 16'h75F0, 16'h5F15, 16'hDFE7, 16'hAE1D,
 16'hAEDE, 16'hC128, 16'hE3D2, 16'hF633,
 16'h1DC8, 16'h753D, 16'h5FBE, 16'hDD48,
 16'hB1B1, 16'hB755, 16'hC0A7, 16'hE95D,
 16'hF99E, 16'h1E66, 16'h7795, 16'h5C71,
 16'hE28A, 16'hB37B, 16'hB67F, 16'hC385,
 16'hE879, 16'hFD88, 16'h1B78, 16'h7388,
 16'h6377, 16'hEC8B, 16'hB673, 16'hB28F,
 16'hC56F, 16'hE492, 16'hF96E, 16'h1992,
 16'h666E, 16'h7192, 16'hFF6E, 16'hB692,
 16'hB66E, 16'hC092, 16'hE16D, 16'hF794,
 16'h0F6C, 16'h5794, 16'h7E6B, 16'h1896,
 16'hBA68, 16'hB69A, 16'hBD65, 16'hDB9D,
 16'hF560, 16'h08A3, 16'h415B, 16'h7FA6,
 16'h345A, 16'hC0A6, 16'hB259, 16'hBEA9,
 16'hD455, 16'hECAD, 16'hFD52, 16'h2BAE,
 16'h7E52, 16'h59AE, 16'hDD53, 16'hB8AC,
 16'hB955, 16'hC6A9, 16'hEB5A, 16'hF9A3,
 16'h1760, 16'h619C, 16'h7369, 16'h0C92,
 16'hB774, 16'hB385, 16'hC281, 16'hDD7A,
 16'hF58B, 16'h0770, 16'h3A95, 16'h7F66,
 16'h3E9F, 16'hCA5C, 16'hB3A8, 16'hBA54,
 16'hD1B0, 16'hEC4D, 16'hFDB6, 16'h1947,
 16'h64BB, 16'h7543, 16'h01C0, 16'hB83D,
 16'hB8C5, 16'hC33A, 16'hDEC7, 16'hF639,
 16'h03C6, 16'h363A, 16'h7EC7, 16'h4438,
 16'hCCC9, 16'hB537, 16'hBBC8, 16'hCE39,
 16'hE8C6, 16'hFD3B, 16'h14C4, 16'h563D,
 16'h7DC1, 16'h1942, 16'hBBBC, 16'hB545,
 16'hBEB9, 16'hD749, 16'hF3B5, 16'hFE4E,
 16'h24AF, 16'h7253, 16'h60AB, 16'hF056,
 16'hB8A9, 16'hB25A, 16'hC1A3, 16'hE05F,
 16'hF69E, 16'h0864, 16'h339C, 16'h7F64,
 16'h499D, 16'hCE60, 16'hB5A3, 16'hB659,
 16'hC6AC, 16'hE54F, 16'hF9B7, 16'h0D41,
 16'h42C7, 16'h7E31, 16'h34D9, 16'hC31D,
 16'hB4EC, 16'hBB0A, 16'hCE00, 16'hEBF7,
 16'hFC13, 16'h0FE2, 16'h4629, 16'h7DCD,
 16'h2B3B, 16'hC1BF, 16'hB247, 16'hB7B3,
 16'hD454, 16'hEBA5, 16'hFD5F, 16'h0FA0,
 16'h4960, 16'h7EA1, 16'h285E, 16'hC0A3,
 16'hB15B, 16'hB9A8, 16'hD453, 16'hEFB4,
 16'hFF46, 16'h11C0, 16'h4539, 16'h7BCE,
 16'h2D2A, 16'hC2E0, 16'hB216, 16'hB8F4,
 16'hD103, 16'hE904, 16'hFAF6, 16'h0A10,
 16'h3DEB, 16'h7C1A, 16'h38E0, 16'hC725,
 16'hB1D7, 16'hB92D, 16'hCECF, 16'hEC34,
 16'hFCCA, 16'h0937, 16'h2FC9, 16'h7836,
 16'h4ECB, 16'hDB35, 16'hB9CB, 16'hBB34,
 16'hC7CD, 16'hE332, 16'hF5D0, 16'h052E,
 16'h1FD4, 16'h6528, 16'h6ADD, 16'h011E,
 16'hB9E7, 16'hB314, 16'hC1F0, 16'hDE0C,
 16'hEFF9, 16'hFE02, 16'h1203, 16'h45F7,
 16'h7B0F, 16'h2DEB, 16'hC21B, 16'hB1E0,
 16'hBC26, 16'hD3D4, 16'hE931, 16'hFFC9,
 16'h083E, 16'h23BC, 16'h734A, 16'h5AB0,
 16'hE756, 16'hB8A3, 16'hB564, 16'hC195,
 16'hE071, 16'hF28B, 16'h0278, 16'h1086,
 16'h467B, 16'h7785, 16'h2A7A, 16'hC287,
 16'hB179, 16'hBC88, 16'hCE76, 16'hEE8C,
 16'hFD71, 16'h0493, 16'h2268, 16'h669E,
 16'h645B, 16'hFCAD, 16'hBA4B, 16'hB0BC,
 16'hC03C, 16'hDDCE, 16'hF028, 16'hFFE2,
 16'h0C13, 16'h30F6, 16'h7802, 16'h4A07,
 16'hDBF0, 16'hBA19, 16'hB4DE, 16'hC82A,
 16'hE2CF, 16'hF537, 16'h03C4, 16'h1241,
 16'h3DBB, 16'h7846, 16'h3ABB, 16'hCA44,
 16'hB4BE, 16'hB83E, 16'hD0C6, 16'hE935,
 16'hF5D2, 16'h0427, 16'h0FE0, 16'h4718,
 16'h7EF1, 16'h3005, 16'hC206, 16'hB5EF,
 16'hBC1B, 16'hCFDC, 16'hED2C, 16'hFACE,
 16'h0838, 16'h0EC1, 16'h4445, 16'h7BB7,
 16'h2C4D, 16'hC6B0, 16'hB551, 16'hBAAF,
 16'hD151, 16'hE9B1, 16'hF64B, 16'h08BA,
 16'h0F40, 16'h3DC7, 16'h7A33, 16'h3AD3,
 16'hCD26, 16'hB4E1, 16'hBF18, 16'hCBF0,
 16'hE608, 16'hF5FE, 16'h04FC, 16'h0F0A,
 16'h30F2, 16'h6F10, 16'h49EF, 16'hE210,
 16'hB5F3, 16'hB50A, 16'hC9FA, 16'hE201,
 16'hF604, 16'h02F8, 16'h090C, 16'h22EF,
 16'h6018, 16'h66DF, 16'h042A, 16'hBBCE,
 16'hB038, 16'hBEC4, 16'hDE3F, 16'hF1BF,
 16'hFE42, 16'h0BBE, 16'h1840, 16'h42C3,
 16'h783A, 16'h31CB, 16'hC72E, 16'hB6DA,
 16'hB61B, 16'hCDF2, 16'hEC01, 16'hF70C,
 16'h05E7, 16'h1026, 16'h26CD, 16'h6140,
 16'h62B3, 16'h015A, 16'hBD9A, 16'hB271,
 16'hBD86, 16'hDB82, 16'hEF78, 16'h008C,
 16'h0A71, 16'h1090, 16'h3B71, 16'h6F8D,
 16'h4676, 16'hDC85, 16'hBA81, 16'hB978,
 16'hC591, 16'hE564, 16'hF5A7, 16'h054E,
 16'h0DBD, 16'h1539, 16'h44D1, 16'h7825,
 16'h33E4, 16'hC714, 16'hB4F3, 16'hB807,
 16'hC5FE, 16'hE4FF, 16'hF002, 16'h00FF,
 16'h06FD, 16'h1009, 16'h43F1, 16'h6D16,
 16'h26E2, 16'hC326, 16'hB1D1, 16'hB73A,
 16'hCBBA, 16'hE651, 16'hF4A4, 16'h0566,
 16'h0B91, 16'h1578, 16'h447F, 16'h7089,
 16'h2970, 16'hC696, 16'hB765, 16'hBC9F,
 16'hD05F, 16'hE6A1, 16'hF361, 16'h039D,
 16'h0D65, 16'h0E99, 16'h3D68, 16'h6F96,
 16'h3A6E, 16'hD78E, 16'hB377, 16'hB983,
 16'hC682, 16'hE37A, 16'hF48A, 16'h0472,
 16'h0D92, 16'h0E6B, 16'h2C96, 16'h646B,
 16'h5393, 16'hF76F, 16'hBB90, 16'hB270,
 16'hC290, 16'hDB71, 16'hF18D, 16'hFE75,
 16'h0689, 16'h0C79, 16'h1B86, 16'h467B,
 16'h6E83, 16'h287F, 16'hC680, 16'hB781,
 16'hB980, 16'hCF7D, 16'hE986, 16'hF777,
 16'h048D, 16'h0A6F, 16'h0E95, 16'h2766,
 16'h5F9F, 16'h595C, 16'h03A9, 16'hBB53,
 16'hAEB1, 16'hC34B, 16'hD9B9, 16'hF042,
 16'hFCC4, 16'h0537, 16'h0ECC, 16'h1231,
 16'h2FD2, 16'h672B, 16'h4BD8, 16'hEB25,
 16'hB5DE, 16'hB320, 16'hC5E1, 16'hDE1D,
 16'hF0E6, 16'hFD18, 16'h0AEA, 16'h1014,
 16'h0FED, 16'h3511, 16'h67F3, 16'h4309,
 16'hE5FA, 16'hB903, 16'hB400, 16'hC6FD,
 16'hDF06, 16'hEEF6, 16'h010F, 16'h0AED,
 16'h0C16, 16'h0DE6, 16'h2E1E, 16'h60DF,
 16'h4C25, 16'hF1D6, 16'hB92E, 16'hB2CF,
 16'hC633, 16'hDDCC, 16'hEF34, 16'hFCCD,
 16'h0732, 16'h0DCE, 16'h0F31, 16'h23D2,
 16'h502B, 16'h5FD9, 16'h1122, 16'hBFE2,
 16'hB31A, 16'hBAEB, 16'hCF0F, 16'hEAF7,
 16'hFB03, 16'h0404, 16'h0BF5, 16'h0B11,
 16'h15E8, 16'h371F, 16'h64DB, 16'h3A2B,
 16'hD8CF, 16'hB636, 16'hB4C6, 16'hC83D,
 16'hDFC0, 16'hF342, 16'h00BD, 16'h0A43,
 16'h08BF, 16'h0D3E, 16'h1FC4, 16'h4539,
 16'h64CC, 16'h1B2F, 16'hC3D7, 16'hB321,
 16'hB5E7, 16'hCE10, 16'hE8FA, 16'hF5FC,
 16'h020E, 16'h06E8, 16'h0C21, 16'h10D7,
 16'h2130, 16'h4BC9, 16'h5C3F, 16'h14B9,
 16'hBF4E, 16'hB2AD, 16'hBE57, 16'hCEA5,
 16'hE85E, 16'hF7A0, 16'h0062, 16'h0B9E,
 16'h0D60, 16'h0AA1, 16'h205F, 16'h48A2,
 16'h5D5D, 16'h1BA5, 16'hBF58, 16'hB4AB,
 16'hBB52, 16'hCAB1, 16'hE64D, 16'hF6B5,
 16'h0249, 16'h0AB8, 16'h1047, 16'h0EBA,
 16'h1A46, 16'h3AB9, 16'h6049, 16'h30B5,
 16'hD94E, 16'hB5AF, 16'hB652, 16'hC5AE,
 16'hDE53, 16'hF3AC, 16'hFC55, 16'h08A9,
 16'h0E58, 16'h0DA9, 16'h0D55, 16'h23AE,
 16'h4B4E, 16'h57B7, 16'h0F43, 16'hBEC5,
 16'hB331, 16'hBDD9, 16'hD41D, 16'hE4EE,
 16'hF608, 16'h0201, 16'h06F5, 16'h0C16,
 16'h0DDE, 16'h132F, 16'h2AC4, 16'h5549,
 16'h45AB, 16'hF960, 16'hBB95, 16'hAF75,
 16'hC083, 16'hD785, 16'hEF75, 16'hF68E,
 16'h026F, 16'h0B94, 16'h096B, 16'h0B95,
 16'h0E6C, 16'h2791, 16'h5074, 16'h4986,
 16'hFF80, 16'hBC79, 16'hB090, 16'hC167,
 16'hD5A3, 16'hE952, 16'hF6B9, 16'h043D,
 16'h0ACC, 16'h0A2D, 16'h0ED9, 16'h0E21,
 16'h1FE5, 16'h4515, 16'h53F1, 16'h1709,
 16'hC5FC, 16'hB501, 16'hBC01, 16'hCDFE,
 16'hE500, 16'hF503, 16'h01FA, 16'h090B,
 16'h07EF, 16'h0916, 16'h0CE4, 16'h1223,
 16'h2CD6, 16'h5031, 16'h40C7, 16'hF442,
 16'hB7B5, 16'hB354, 16'hC6A3, 16'hD865,
 16'hEE94, 16'hFA72, 16'hFF89, 16'h087B,
 16'h0B82, 16'h0F81, 16'h117C, 16'h1287,
 16'h3076, 16'h538C, 16'h3773, 16'hEC8E,
 16'hB873, 16'hB28B, 16'hC576, 16'hDC89,
 16'hED79, 16'hFB85, 16'h077E, 16'h087F,
 16'h0884, 16'h0E79, 16'h0E89, 16'h1275,
 16'h2A8D, 16'h4973, 16'h458C, 16'hFF75,
 16'hBC8A, 16'hB276, 16'hBE8B, 16'hD475,
 16'hEB8A, 16'hF878, 16'h0385, 16'h0A7E,
 16'h0B7F, 16'h0E84, 16'h0E78, 16'h0C8C,
 16'h1671, 16'h3890, 16'h4F70, 16'h228F,
 16'hD873, 16'hB58A, 16'hB57A, 16'hCA81,
 16'hDE85, 16'hF075, 16'hFF91, 16'h0368,
 16'h0BA0, 16'h0A58, 16'h0EB1, 16'h0D45,
 16'h0BC5, 16'h1D31, 16'h36D9, 16'h4D1E,
 16'h1DEA, 16'hD40E, 16'hB9F9, 16'hB402,
 16'hC802, 16'hE1FB, 16'hF307, 16'h00F7,
 16'h0A09, 16'h0EF9, 16'h0E04, 16'h1101,
 16'h0BF8, 16'h0810, 16'h12E7, 16'h3023,
 16'h47D3, 16'h3437, 16'hEEBF, 16'hB84B,
 16'hB2AB, 16'hC55F, 16'hDB98, 16'hEE6F,
 16'hFC8B, 16'h0379, 16'h0B86, 16'h0E79,
 16'h0E89, 16'h0E72, 16'h0A96, 16'h0B60,
 16'h19AD, 16'h3644, 16'h4CCB, 16'h1C25,
 16'hD3EC, 16'hB602, 16'hB211, 16'hC5DC,
 16'hDB38, 16'hE9B3, 16'hFC61, 16'h048C,
 16'h0786, 16'h0D6B, 16'h0BA2, 16'h0852,
 16'h07B7, 16'h0644, 16'h0FBE, 16'h3342,
 16'h47BC, 16'h2248, 16'hE2B3, 16'hB654,
 16'hB1A1, 16'hCA6D, 16'hD984, 16'hEE8D,
 16'hFD61, 16'h03B0, 16'h0B3F, 16'h0AD2,
 16'h0F1E, 16'h0BF2, 16'h09FE, 16'h0911,
 16'h06E2, 16'h1C29, 16'h3BCF, 16'h4237,
 16'h0FC5, 16'hCB3D, 16'hB5C2, 16'hB73E,
 16'hCFC6, 16'hE333, 16'hF1D4, 16'h0424,
 16'h08E5, 16'h0E12, 16'h0DF8, 16'h0CFD,
 16'h0B0E, 16'h0BE7, 16'h0823, 16'h06D4,
 16'h1934, 16'h36C6, 16'h453F, 16'h18BD,
 16'hD445, 16'hB8BA, 16'hB746, 16'hCCBC,
 16'hE141, 16'hF2C3, 16'hFF38, 16'h08CE,
 16'h0E2B, 16'h0ADC, 16'h101C, 16'h09ED,
 16'h080A, 16'h08FE, 16'h0AFB, 16'h0E0C,
 16'h20EE, 16'h3917, 16'h37E4, 16'h0B20,
 16'hC8DE, 16'hB624, 16'hBEDB, 16'hCF24,
 16'hE4DF, 16'hF41B, 16'hFFED, 16'h0B0B,
 16'h0AFD, 16'h0AFA, 16'h100F, 16'h0AE8,
 16'h0B22, 16'h07D4, 16'h0635, 16'h07C3,
 16'h1544, 16'h2FB5, 16'h4052, 16'h20A7,
 16'hDF60, 16'hB99B, 16'hB467, 16'hCC98,
 16'hE068, 16'hF199, 16'hFB66, 16'h029C,
 16'h0E60, 16'h0AA6, 16'h0B52, 16'h0DB7,
 16'h0D3F, 16'h06CC, 16'h0929, 16'h06E2,
 16'h0111, 16'h15FD, 16'h2FF5, 16'h3C18,
 16'h1EDC, 16'hE42F, 16'hB9C6, 16'hB546,
 16'hC7AE, 16'hDB5C, 16'hED9D, 16'hFA69,
 16'h0591, 16'h0975, 16'h0D86, 16'h0E7E,
 16'h0D7F, 16'h0A83, 16'h077C, 16'h0884,
 16'h057E, 16'h027E, 16'h0386, 16'h1977,
 16'h2E8C, 16'h3870, 16'h1495, 16'hD666,
 16'hBC9E, 16'hB65F, 16'hCCA3, 16'hDE5B,
 16'hEFA8, 16'h0054, 16'h06B0, 16'h0A4D,
 16'h09B5, 16'h0E4A, 16'h0AB6, 16'h0B4B,
 16'h07B4, 16'h094C, 16'h06B4, 16'h044C,
 16'hFEB4, 16'h094E, 16'h20AE, 16'h3155,
 16'h36A8, 16'h035C, 16'hCAA1, 16'hB462,
 16'hBB9A, 16'hD06A, 16'hE492, 16'hF573,
 16'h0187, 16'h0780, 16'h0B79, 16'h0A8E,
 16'h0E6A, 16'h0B9F, 16'h0657, 16'h08B4,
 16'h0741, 16'h02C9, 16'hFF2E, 16'h04DC,
 16'hFE19, 16'h0CF2, 16'h2602, 16'h350A,
 16'h25EB, 16'hF320, 16'hC4D6, 16'hB631,
 16'hC1C9, 16'hD53C, 16'hEAC1, 16'hF741,
 16'h06BD, 16'h0843, 16'h0CC0, 16'h0E3C,
 16'h09CA, 16'h0E2D, 16'h0ADE, 16'h0416,
 16'h05F7, 16'h04FC, 16'h0111, 16'h01E2,
 16'hFD2B, 16'h00C7, 16'h1149, 16'h28A6,
 16'h356B, 16'h1C85, 16'hE889, 16'hC46B,
 16'hB7A0, 16'hC156, 16'hDAB3, 16'hEA46,
 16'hFABE, 16'h0440, 16'h07C1, 16'h0D3F,
 16'h0BC1, 16'h0B40, 16'h08BE, 16'h0A45,
 16'h04B8, 16'h004C, 16'h04AF, 16'h0256,
 16'hFCA5, 16'h0160, 16'h019D, 16'hFD65,
 16'h1199, 16'h2669, 16'h2F95, 16'h1F6C,
 16'hF095, 16'hC668, 16'hB69D, 16'hC05E,
 16'hD6A8, 16'hE850, 16'hF6B9, 16'h043E,
 16'h0ACB, 16'h0C2D, 16'h0BDA, 16'h081F,
 16'h0BE9, 16'h0A0D, 16'h01FD, 16'h03F9,
 16'h0110, 16'h00E9, 16'h031C, 16'h03E0,
 16'h0023, 16'hFDDA, 16'h0129, 16'h0AD5,
 16'h192C, 16'h26D5, 16'h2D29, 16'h0DDA,
 16'hDE22, 16'hC2E3, 16'hB918, 16'hC7EE,
 16'hDF0B, 16'hEEFD, 16'hFCFB, 16'h040C,
 16'h0AED, 16'h0E19, 16'h0AE2, 16'h0C24,
 16'h0AD4, 16'h0834, 16'h07C5, 16'h0242,
 16'h05B7, 16'h044E, 16'hFEAD, 16'h0059,
 16'hFEA2, 16'hFE63, 16'h0197, 16'hFD6F,
 16'h038B, 16'h167A, 16'h2182, 16'h2D82,
 16'h1F7C, 16'hF685, 16'hCE79, 16'hBB89,
 16'hC276, 16'hD38C, 16'hE573, 16'hF78D,
 16'h0073, 16'h068C, 16'h0B77, 16'h0B85,
 16'h0D80, 16'h0D7B, 16'h0B8A, 16'h0371,
 16'h0694, 16'h0166, 16'h01A0, 16'h045B,
 16'h00AB, 16'hFF4E, 16'hFDBA, 16'h023D,
 16'h00CC, 16'hFE2C, 16'hFBDC, 16'h021C,
 16'h08EC, 16'h1B0C, 16'h22FC, 16'h28FB,
 16'h120D, 16'hE4EC, 16'hCA1B, 16'hB9DF,
 16'hC826, 16'hD7D4, 16'hED32, 16'hF8C9,
 16'h023B, 16'h09C3, 16'h0C3E, 16'h0BC2,
 16'h0A3D, 16'h08C5, 16'h0738, 16'h08CC,
 16'h012F, 16'h06D7, 16'h0322, 16'hFFE6,
 16'h0111, 16'hFFF9, 16'h03FC, 16'h0010,
 16'hFDE3, 16'hFF2A, 16'hFCCA, 16'h0141,
 16'h01B4, 16'hFF58, 16'h069B, 16'h1571,
 16'h1E84, 16'h2385, 16'h2275, 16'hFD8F,
 16'hD96F, 16'hC191, 16'hBD70, 16'hCB8E,
 16'hDD77, 16'hF381, 16'hFA88, 16'h046E,
 16'h0A9E, 16'h0E55, 16'h0DB9, 16'h0C37,
 16'h0ADB, 16'h0112, 16'h0401, 16'hFFEC,
 16'h0027, 16'hFFC6, 16'hFA4D, 16'h00A1,
 16'h006F, 16'hFC83, 16'hFA89, 16'hFD6D,
 16'hFE9B, 16'hFC5E, 16'hFDA8, 16'h0055,
 16'hFCAB, 16'hFC58, 16'hFCA2, 16'hFD66,
 16'h0691, 16'h0E79, 16'h197C, 16'h1E91,
 16'h1C5F, 16'h06B2, 16'hE53D, 16'hCDD4,
 16'hBC1A, 16'hC6F9, 16'hD8F3, 16'hE921,
 16'hF7CB, 16'h0048, 16'h08A7, 16'h0A69,
 16'h0E88, 16'h0D84, 16'h0D73, 16'h0B95,
 16'h0A64, 16'h08A2, 16'h0259, 16'h00AA,
 16'h0357, 16'h00A5, 16'hFE61, 16'h0498,
 16'hFE70, 16'hFE87, 16'h0384, 16'hFD70,
 16'hFD9C, 16'h0158, 16'hFFB3, 16'hFD43,
 16'hFDC7, 16'hFE2F, 16'hFFDA, 16'h001E,
 16'hFFE9, 16'hFD12, 16'h00F2, 16'h020A,
 16'h0AF8, 16'h1808, 16'h17F6, 16'h1C0E,
 16'h15ED, 16'hFE19, 16'hE2E0, 16'hD228,
 16'hC0CE, 16'hC53C, 16'hD8BB, 16'hE94D,
 16'hF7AC, 16'h045B, 16'h0A9E, 16'h0C68,
 16'h0E92, 16'h0C73, 16'h0A8A, 16'h0977,
 16'h098A, 16'h0473, 16'h0791, 16'h046B,
 16'h009A, 16'hFF5F, 16'h04A9, 16'h014E,
 16'hFFBD, 16'h0338, 16'hFFD2, 16'hFD24,
 16'hFCE5, 16'h0113, 16'hFEF4, 16'h0406,
 16'hFF00, 16'hFDF9, 16'h010D, 16'hFDEF,
 16'hFD14, 16'hFDEB, 16'hFC14, 16'hFCED,
 16'hFC13, 16'hFDEE, 16'h0010, 16'hFFF3,
 16'h0008, 16'hFFFE, 16'hFFFC, 16'h000A,
 16'h0DF1, 16'h0F13, 16'h14E9, 16'h131A,
 16'h0EE4, 16'h051E, 16'hEAE1, 16'hDB20,
 16'hCDDF, 16'hC621, 16'hCCE0, 16'hE01D,
 16'hE9E7, 16'hFB15, 16'h04EF, 16'h0B0D,
 16'h0FF6, 16'h0B06, 16'h0C00, 16'h09FA,
 16'h090B, 16'h0AF0, 16'h0314, 16'h18EA,
 16'h2F18, 16'hF6E6, 16'hE51B, 16'hF0E5,
 16'hF01A, 16'hF3E8, 16'h0115, 16'h25EF,
 16'hFA0C, 16'hE1FA, 16'h01FE, 16'hF00B,
 16'h03EB, 16'h2621, 16'hF5D3, 16'hE639,
 16'h01BA, 16'hEE53, 16'h07A1, 16'h256B,
 16'hF28B, 16'hE87E, 16'h007A, 16'hEF8C,
 16'h026F, 16'h2094, 16'hF76C, 16'hE592,
 16'hFF72, 16'hF388, 16'h007F, 16'h2078,
 16'hF694, 16'hE55E, 16'hFFB3, 16'hED39,
 16'h00DC, 16'h230E, 16'hF70B, 16'hE7DB,
 16'h0040, 16'hEBA4, 16'h0277, 16'h236F,
 16'hF3AB, 16'hE43C, 16'h00DC, 16'hEE0E,
 16'h0205, 16'h22EA, 16'hF425, 16'hEACF,
 16'h013A, 16'hEDBF, 16'h0046, 16'h1DB8,
 16'hF747, 16'hEEBC, 16'h013F, 16'hEDC9,
 16'hFD2C, 16'h1BE0, 16'hF911, 16'hF302,
 16'hFFEA, 16'hE92A, 16'hFDC1, 16'h1554,
 16'h0297, 16'hFA7F, 16'hF86A, 16'hEEAD,
 16'hF83D, 16'h0AD8, 16'h1214, 16'hFDFF,
 16'hF0EE, 16'hF324, 16'hF6CC, 16'h0442,
 16'h18B1, 16'hFE5A, 16'hE89C, 16'hF86D,
 16'hEF8B, 16'h047C, 16'h1E7E, 16'hFA86,
 16'hE477, 16'h008A, 16'hEB78, 16'hFE85,
 16'h227F, 16'hF37B, 16'hED8C, 16'h016B,
 16'hEC9F, 16'hFD57, 16'h19B4, 16'hFC41,
 16'hF6C9, 16'hFA2D, 16'hEEDE, 16'hF717,
 16'h0AF4, 16'h1101, 16'hFE0A, 16'hECED,
 16'hF71A, 16'hF3E0, 16'h0425, 16'h22D8,
 16'hF629, 16'hE4D7, 16'h0027, 16'hEBDE,
 16'hFD1C, 16'h22EA, 16'hF60E, 16'hEBFB,
 16'hFFFB, 16'hEE11, 16'hFCE3, 16'h1428,
 16'h01CD, 16'hFA3E, 16'hF5B7, 16'hF354,
 16'hF9A2, 16'h0367, 16'h1E92, 16'h0073,
 16'hEA8A, 16'hFD76, 16'hED8D, 16'h046F,
 16'h2396, 16'hF564, 16'hECA3, 16'h0154,
 16'hEDB7, 16'hFD3D, 16'h15CF, 16'h0325,
 16'hFFE7, 16'hF60D, 16'hEFFE, 16'hF5F9,
 16'h040F, 16'h1DEA, 16'hFB1B, 16'hE8E1,
 16'h0022, 16'hEEDD, 16'h0022, 16'h1EE1,
 16'hF719, 16'hF5EF, 16'hFC08, 16'hF001,
 16'hF9F7, 16'h0A12, 16'h15E3, 16'hFE28,
 16'hEDCD, 16'hFD3E, 16'hF1B9, 16'h014E,
 16'h22AC, 16'hF459, 16'hEFA3, 16'hFF5F,
 16'hEEA2, 16'hFC5B, 16'h0FAA, 16'h0D4F,
 16'hFFB9, 16'hF03E, 16'hF5CD, 16'hF326,
 16'h01E9, 16'h2306, 16'hF80C, 16'hE9E2,
 16'hFD30, 16'hF2BF, 16'hFD51, 16'h11A0,
 16'h0A6F, 16'hFA82, 16'hF08C, 16'hF968,
 16'hF3A2, 16'h0156, 16'h25AF, 16'hF54E,
 16'hE9B4, 16'h004C, 16'hF0B1, 16'hFB53,
 16'h10A8, 16'h0D5F, 16'h0199, 16'hF370,
 16'hF685, 16'hF588, 16'h016A, 16'h1FA4,
 16'hF34E, 16'hF3BF, 16'hFD35, 16'hF2D7,
 16'hFE1E, 16'h03EB, 16'h1A0C, 16'hFEFD,
 16'hECFC, 16'hFD09, 16'hF3F2, 16'hFF12,
 16'h18EB, 16'hFD18, 16'hF7E6, 16'hF71A,
 16'hF5E7, 16'hF716, 16'h03ED, 16'h2610,
 16'hF8F5, 16'hED06, 16'hFCFD, 16'hF000,
 16'hF702, 16'h07FE, 16'h0B02, 16'hFBFE,
 16'hED01, 16'hF301, 16'hF4FD, 16'hFB07,
 16'h18F3, 16'hFA13, 16'hF3E7, 16'hF721,
 16'hEFD6, 16'hF933, 16'h00C3, 16'h2247,
 16'hF6B1, 16'hEB56, 16'hFAA3, 16'hF063,
 16'hFB99, 16'h0869, 16'h1697, 16'hFE67,
 16'hEF9D, 16'hFA5E, 16'hF4A8, 16'hFA50,
 16'h14BA, 16'h0439, 16'hFBD8, 16'hF715,
 16'hF2FF, 16'hF3EB, 16'h022B, 16'h1BC1,
 16'hF754, 16'hF596, 16'hFA80, 16'hF56A,
 16'hF9AB, 16'h0343, 16'h1FCD, 16'hF725,
 16'hECE7, 16'hFC0F, 16'hF2F8, 16'hFC04,
 16'h08FF, 16'h1B00, 16'hFAFD, 16'hEE0A,
 16'hFAEC, 16'hF521, 16'hFDD1, 16'h0A3E,
 16'h0DB1, 16'hFF61, 16'hF38B, 16'hF68B,
 16'hF55F, 16'hFFB8, 16'h1230, 16'h03E7,
 16'hF904, 16'hF310, 16'hF5DE, 16'hFA31,
 16'hFFC3, 16'h1748, 16'hFFAF, 16'hF757,
 16'hFCA4, 16'hF360, 16'hF39F, 16'h0360,
 16'h18A2, 16'hF75A, 16'hF7AD, 16'hFA4A,
 16'hF5C0, 16'hF936, 16'hFFD5, 16'h1C1F,
 16'hF9ED, 16'hF708, 16'hFC02, 16'hF6F4,
 16'hFA16, 16'h00E0, 16'h1E29, 16'hF3CF,
 16'hF337, 16'hFDC5, 16'hF63E, 16'hFAC0,
 16'h0041, 16'h1EBF, 16'hF440, 16'hF2C2,
 16'hFE3C, 16'hF6C7, 16'hF734, 16'h03D3,
 16'h1E26, 16'hF3E0, 16'hF61A, 16'hFCEA,
 16'hF614, 16'hF7ED, 16'h0412, 16'h19EE,
 16'hF612, 16'hF5EE, 16'hFA13, 16'hF9EB,
 16'hFB18, 16'hFFE3, 16'h1924, 16'hF6D4,
 16'hF835, 16'hFAC3, 16'hF544, 16'hF9B5,
 16'h0052, 16'h16A7, 16'hF860, 16'hFC99,
 16'hFC6D, 16'hF38E, 16'hFA76, 16'hFD88,
 16'h1078, 16'h0089, 16'hF875, 16'hF68F,
 16'hF16C, 16'hF899, 16'hFE62, 16'h0EA5,
 16'h0952, 16'hF9B8, 16'hF53C, 16'hF5D1,
 16'hFB23, 16'hF6E9, 16'h070A, 16'h1204,
 16'hFCEC, 16'hF725, 16'hF6CB, 16'hF945,
 16'hF7AC, 16'h0361, 16'h1992, 16'hF97B,
 16'hF27A, 16'hFA90, 16'hF566, 16'hF7A3,
 16'h0256, 16'h1AAF, 16'hF54E, 16'hF1B3,
 16'hFA4D, 16'hF2B4, 16'hFD4B, 16'h03B5,
 16'h114C, 16'hF9B2, 16'hFC52, 16'hFAAA,
 16'hF15A, 16'hFAA0, 16'hFB67, 16'h0992,
 16'h0D76, 16'hFE83, 16'hF682, 16'hF679,
 16'hFC8B, 16'hF773, 16'h038F, 16'h1A70,
 16'hF890, 16'hF371, 16'hFC8C, 16'hFB78,
 16'hF883, 16'h0183, 16'h1777, 16'hFA8F,
 16'hF56A, 16'hFD9D, 16'hF65B, 16'hFAAD,
 16'hFD4B, 16'h0ABD, 16'h0D3C, 16'hFACA,
 16'hF632, 16'hF6CF, 16'hFC32, 16'hF5CC,
 16'h0338, 16'h19C3, 16'hF544, 16'hF5B2,
 16'hFC5A, 16'hF398, 16'hFD7A, 16'hFE72,
 16'h0AA3, 16'h0446, 16'hFBD2, 16'hFB16,
 16'hF404, 16'hFAE1, 16'hF738, 16'h03B1,
 16'h1A65, 16'hF887, 16'hF18D, 16'hF860,
 16'hF6B0, 16'hF843, 16'hFFC7, 16'h1132,
 16'hFDD4, 16'hFA28, 16'hF9D9, 16'hF229,
 16'hFDD1, 16'hF738, 16'h03BC, 16'h1853,
 16'hF39D, 16'hF374, 16'hFA7A, 16'hF596,
 16'hF95B, 16'hFFB4, 16'h0E3F, 16'hFFCC,
 16'hFB29, 16'hFBE0, 16'hF41B, 16'hF9E8,
 16'hF817, 16'h02E7, 16'h191E, 16'hF3DB,
 16'hF42F, 16'hFFC4, 16'hF44B, 16'hFDA6,
 16'hFD6A, 16'h0A83, 16'h0891, 16'hF95A,
 16'hF7BD, 16'hF62C, 16'hF9E9, 16'hF703,
 16'h040F, 16'h13E2, 16'hF82B, 16'hFBCA,
 16'hFD3D, 16'hF2BE, 16'h0145, 16'hF8BB,
 16'h0143, 16'h17C1, 16'hFB37, 16'hF5D5,
 16'hFD1C, 16'hF5F5, 16'hFFF9, 16'hFA1A,
 16'h08D1, 16'h0F47, 16'hFF9E, 16'hF77E,
 16'hF566, 16'hF9B6, 16'hFB2E, 16'hFFEE,
 16'h0DF6, 16'hFE26, 16'hF8C0, 16'hFD59,
 16'hF58F, 16'h0188, 16'hF461, 16'h04B5,
 16'h1337, 16'hF7DB, 16'hF916, 16'hFDF6,
 16'hF600, 16'h0109, 16'hF8EF, 16'h0117,
 16'h17E5, 16'hF91D, 16'hF6E4, 16'hFE19,
 16'hF4EC, 16'h020C, 16'hFDFD, 16'h01F9,
 16'h1412, 16'hFAE4, 16'hF826, 16'hFDCE,
 16'hF63F, 16'h01B4, 16'hFB59, 16'h049B,
 16'h0971, 16'hFA83, 16'hF788, 16'hF76E,
 16'hFC9B, 16'hFD5E, 16'h00A8, 16'h0C52,
 16'h08B5, 16'h0045, 16'hF7BF, 16'hF83D,
 16'hFDC7, 16'hFE37, 16'hFDCB, 16'h0832,
 16'h08D0, 16'hFA2F, 16'hF9D3, 16'hFC2B,
 16'hFCD7, 16'hFD26, 16'h00DE, 16'h061D,
 16'h08E8, 16'hFF14, 16'hF7F0, 16'hF70C,
 16'hFAF8, 16'h0003, 16'h0002, 16'h06FA,
 16'h090A, 16'hFCF2, 16'hF811, 16'hFBEC,
 16'hFC17, 16'hFCE6, 16'hFC1C, 16'h06E3,
 16'h0C1C, 16'hFEE7, 16'hF815, 16'hFCF0,
 16'hFC0A, 16'hFCFC, 16'hFCFE, 16'h0409,
 16'h0FF0, 16'hFF17, 16'hF2E1, 16'hF727,
 16'hF2D1, 16'hFA37, 16'hFAC2, 16'h0044,
 16'h0FB6, 16'hF54F, 16'hF2AE, 16'hFC54,
 16'hF5AB, 16'hFE53, 16'hF6B1, 16'h024A,
 16'h0FBD, 16'hF53A, 16'hF9D0, 16'h0025,
 16'hF2E8, 16'h0009, 16'hF908, 16'h00E5,
 16'h0B31, 16'hF7B7, 16'hFD62, 16'hFC85,
 16'hF695, 16'hFF51, 16'hFBC9, 16'h001D,
 16'h07FC, 16'h02EE, 16'hFD27, 16'hFBC4,
 16'hFB4E, 16'hF8A2, 16'h016C, 16'hFD89,
 16'h027F, 16'h0C7B, 16'hFC88, 16'hF779,
 16'hFE81, 16'hF989, 16'h006C, 16'hFBA1,
 16'hFD4F, 16'h0CC3, 16'hF828, 16'hFBF0,
 16'hFCF7, 16'hFA22, 16'hFFC3, 16'hFF58,
 16'h008D, 16'h038E, 16'h0759, 16'hFDBD,
 16'hF92F, 16'hFCE4, 16'hFA0B, 16'h0003,
 16'hFBF2, 16'h0116, 16'h0EE6, 16'hF61B,
 16'hFBE5, 16'hFD19, 16'hF9EB, 16'h0010,
 16'hFFF6, 16'h0002, 16'h0307, 16'h07EF,
 16'hFD1A, 16'hF8DF, 16'hFD27, 16'hF9D4,
 16'h0030, 16'hFECC, 16'h0137, 16'h0DC8,
 16'hF739, 16'hFCC7, 16'hFC37, 16'hFACD,
 16'hFF2D, 16'hFFDA, 16'hFF1F, 16'h00E9,
 16'h080F, 16'hFDF8, 16'hFA01, 16'hFC05,
 16'hFCF6, 16'hFC0F, 16'hFDEE, 16'h0112,
 16'h0CF0, 16'hFA0B, 16'hFCFC, 16'hFCFD,
 16'hFA0B, 16'hFFEB, 16'hFD21, 16'hFED0,
 16'h0141, 16'h0CAF, 16'hF761, 16'hF98E,
 16'hFD82, 16'hFA6F, 16'hFBA1, 16'hFF51,
 16'hFFBA, 16'h003C, 16'h08CC, 16'hFC2E,
 16'hFCD6, 16'hFC29, 16'hFAD6, 16'hFF2D,
 16'hFFCD, 16'hFF3B, 16'h04BC, 16'h014E,
 16'hFAA7, 16'hFC65, 16'hFC8E, 16'hFC80,
 16'hFD71, 16'hFD9E, 16'hFD54, 16'h07B9,
 16'hFD3A, 16'hFCD1, 16'hFC26, 16'hFAE2,
 16'hFB17, 16'hFEEE, 16'h000F, 16'hFEF1,
 16'h0912, 16'hF6E9, 16'hFB1D, 16'hF9DD,
 16'hFB29, 16'hFCD0, 16'h0039, 16'hFFBD,
 16'hFF4E, 16'h08A7, 16'hF863, 16'hFB93,
 16'hFD76, 16'hFB83, 16'hFB84, 16'hFF77,
 16'hFF8A, 16'hFF77, 16'h0787, 16'hFA7D,
 16'hFA7E, 16'hFF86, 16'hF677, 16'hFC8D,
 16'h006E, 16'hFE98, 16'h005F, 16'h06AC,
 16'hFB4A, 16'hF9C0, 16'h0036, 16'hF9D3,
 16'hFB25, 16'hFAE2, 16'hFA19, 16'h00EB,
 16'h0811, 16'hF9F2, 16'hFD0C, 16'hFBF4,
 16'hF70E, 16'hFFEF, 16'h0015, 16'hF9E5,
 16'h0220, 16'h06DB, 16'h012B, 16'h01CF,
 16'hF836, 16'hFBC5, 16'hFD40, 16'hFBBA,
 16'hFD4D, 16'hFBAC, 16'h015B, 16'h05A0,
 16'hFD63, 16'hFC9A, 16'hFD69, 16'hFC94,
 16'hFA6E, 16'hFF92, 16'hFF6E, 16'hFF91,
 16'h086F, 16'hF792, 16'hFA6D, 16'hFF95,
 16'hFC69, 16'hFF99, 16'h0064, 16'hFBA1,
 16'hFD59, 16'h02AE, 16'hFD4A, 16'hFBBD,
 16'hFD3D, 16'hFCC9, 16'hFD31, 16'hFDD5,
 16'hFE23, 16'hFCE6, 16'hFE11, 16'h07F8,
 16'hFCFF, 16'hF80A, 16'hFCEC, 16'hFD1F,
 16'hFAD5, 16'hFF37, 16'hFFBF, 16'hFF48,
 16'h07B2, 16'hFA54, 16'hFCA7, 16'hFC5D,
 16'hFAA1, 16'hFF5E, 16'hFAA5, 16'h0057,
 16'hFEAF, 16'h004A, 16'h03BF, 16'hFE35,
 16'hFBD9, 16'hFD18, 16'hFBF9, 16'hFAF5,
 16'hFF1D, 16'hFAD1, 16'hFF42, 16'h04AB,
 16'hFA67, 16'hFC87, 16'hFD8A, 16'hF967,
 16'h00A8, 16'hFF4A, 16'hFFC2, 16'hFF32,
 16'h00D9, 16'h061F, 16'hFAE7, 16'hFC15,
 16'hFCED, 16'hFC12, 16'hFCED, 16'hFD16,
 16'hFDE5, 16'hFD21, 16'h02D9, 16'h052E,
 16'hFDC8, 16'hFB44, 16'hFDAE, 16'hFB61,
 16'hFD91, 16'hFC7C, 16'hFE76, 16'hFD99,
 16'h0159, 16'h01B4, 16'hFC3F, 16'hFCCE,
 16'hFC25, 16'hFCE9, 16'hFD09, 16'hFE04,
 16'hFCEF, 16'hFE1D, 16'h00D8, 16'h0133,
 16'hFBC4, 16'hFD42, 16'hFCB9, 16'hFC4B,
 16'hFDB3, 16'hFD4F, 16'hFDAF, 16'hFD51,
 16'h03B1, 16'hFD4C, 16'hFBB9, 16'hFD41,
 16'hFBC5, 16'hFE33, 16'hFCD6, 16'hFE21,
 16'hFCEA, 16'h0209, 16'h0104, 16'hFAEE,
 16'h0021, 16'hFCD2, 16'hFC3A, 16'h00BA,
 16'hFC52, 16'hFCA2, 16'hFC6A, 16'hFC8C,
 16'h017C, 16'hFF7D, 16'hFD89, 16'hFC72,
 16'hFC92, 16'hFC6D, 16'hFD90, 16'hFD75,
 16'hFD84, 16'h0185, 16'h0172, 16'h0198,
 16'hFD5C, 16'hFCB1, 16'hFC40, 16'hFCD1,
 16'hFD1D, 16'hFCF5, 16'h00F9, 16'hFC1A,
 16'h00D2, 16'h0641, 16'hFCAC, 16'hFD66,
 16'h008B, 16'hFD82, 16'hFC71, 16'hFC9B,
 16'h005B, 16'hFCAD, 16'h004D, 16'h02B8,
 16'hF945, 16'hFDBB, 16'hFF47, 16'hFDB5,
 16'hFF52, 16'hFDA6, 16'hFB62, 16'hFD94,
 16'h0077, 16'h007E, 16'h018D, 16'hFA68,
 16'hFCA2, 16'hFC53, 16'hFCB8, 16'hFD3E,
 16'hFDCB, 16'hFE2D, 16'hF8DA, 16'h0120,
 16'hFFE4, 16'hFA1A, 16'hFAE7, 16'hFA1A,
 16'hF9E4, 16'hFD1E, 16'hF9DD, 16'hFE2B,
 16'hFECC, 16'hFB3E, 16'hFEB7, 16'h0053,
 16'hFEA3, 16'hFB68, 16'hFE8D, 16'hFB7D,
 16'hFE7A, 16'h008E, 16'hFE6C, 16'h009A,
 16'hFE5F, 16'h01A7, 16'h0055, 16'hFCAD,
 16'h0053, 16'hFCAB, 16'hFC59, 16'hFCA2,
 16'hFC64, 16'hFE94, 16'hFC75, 16'hFE82,
 16'h0088, 16'hFD6D, 16'hFC9E, 16'hFC58,
 16'hFDB2, 16'hFE44, 16'hFDC5, 16'hFE33,
 16'hFED4, 16'h0026, 16'hFFE0, 16'h011A,
 16'hFCEB, 16'hFD11, 16'hFCF2, 16'hFC0C,
 16'hFDF4, 16'hFD0D, 16'hFDF1, 16'hFD12,
 16'hFDEB, 16'h0117, 16'h00E6, 16'hFD1E,
 16'hFBDE, 16'hFD25, 16'hFCD9, 16'h0129,
 16'hFCD5, 16'hFC2C, 16'h00D3, 16'hFC2E,
 16'h00D2, 16'h002D, 16'hFCD4, 16'hFD2C,
 16'hFCD4, 16'hFC2C, 16'hFDD4, 16'hFD2B,
 16'hFDD6, 16'h012A, 16'hFCD5, 16'hFC2D,
 16'h00CF, 16'hFC36, 16'hFCC5, 16'hFD40,
 16'hFBBA, 16'h024C, 16'hFBAF, 16'hFD57,
 16'hFBA2, 16'hFD65, 16'h0094, 16'hFD73,
 16'h0086, 16'hFD81, 16'h0078, 16'h018E,
 16'hFC6D, 16'hFD98, 16'hFF64, 16'hFD9E,
 16'hFF61, 16'hFDA0, 16'hFF61, 16'h019C,
 16'hFC68, 16'hFC93, 16'hFC74, 16'hFC84,
 16'h0085, 16'hFC70, 16'hFC9C, 16'hFC58,
 16'hFDB4, 16'hFF40, 16'hFFCC, 16'h0028,
 16'hFCE5, 16'h010D, 16'hFD01, 16'hFCF1

};
assign depth = 4080; // same as numbers of samples
/* end sine 441 hz*/



assign dout[15:0] = ROM[adress][15:0]; // take the adress row
assign repeats = 1; // repeat once
endmodule


