module player_ROM (
	
	input clk,
	input resetN,
	input [31:0] adress, // for future purpose
	output [15:0] dout,
	output [17:0] depth,
	output [31:0] repeats

);
/* player_explosion sound*/
 // stroe the value
bit [0:8730][15:0] player_ROM ={ // need to be 0 to 102 so first 2 bytes be on the left 
16'hF9DF, 16'hF6A9, 16'hF714, 16'hF70E,
 16'hF7DC, 16'hF835, 16'h00BC, 16'h0251,
 16'h04A3, 16'h0168, 16'hFC8F, 16'hF779,
 16'hF67E, 16'hF78B, 16'hFC6C, 16'h009D,
 16'h065A, 16'h09AE, 16'h044B, 16'hFBBC,
 16'hEC3D, 16'hE3CB, 16'hDA2C, 16'hDCDC,
 16'hE41D, 16'hF4EA, 16'h0612, 16'h0CF1,
 16'h0E0A, 16'h02FA, 16'hFA03, 16'hEA01,
 16'hDEFC, 16'hDA04, 16'hDAFD, 16'hEA02,
 16'hF200, 16'hF4FC, 16'hF70A, 16'hF7EE,
 16'h011C, 16'h05DA, 16'h0A30, 16'h15C4,
 16'h224A, 16'h2BA8, 16'h2D67, 16'h2D89,
 16'h2086, 16'h0F6B, 16'h04A6, 16'hF349,
 16'hE2C7, 16'hCF28, 16'hC7EA, 16'hCB06,
 16'hCF09, 16'hD1E8, 16'hD725, 16'hE6D0,
 16'hFD3A, 16'h0EBE, 16'h0B48, 16'h08B3,
 16'h0950, 16'h14AE, 16'h2354, 16'h2CAA,
 16'h2858, 16'h18A6, 16'h055B, 16'hEEA6,
 16'hE957, 16'hE9AD, 16'hED50, 16'hF6B2,
 16'h094D, 16'h14B4, 16'h0C4B, 16'h04B5,
 16'h054B, 16'h0EB6, 16'h1A4A, 16'h27B5,
 16'h374B, 16'h3AB4, 16'h3C4E, 16'h37B0,
 16'h2D53, 16'h22AA, 16'h0F58, 16'hF0A4,
 16'hCB61, 16'hA69B, 16'h8569, 16'h8000,
 16'h806E, 16'h8291, 16'h8970, 16'h928F,
 16'hAE72, 16'hD18E, 16'hE971, 16'hF790,
 16'h076F, 16'h0A92, 16'h106D, 16'h2C96,
 16'h4365, 16'h4FA0, 16'h535A, 16'h49AD,
 16'h3F4C, 16'h34BB, 16'h353D, 16'h49CC,
 16'h6C2A, 16'h7EE1, 16'h7F14, 16'h7EF7,
 16'h7EFE, 16'h7F0D, 16'h6FE8, 16'h5423,
 16'h3FD3, 16'h2B35, 16'h01C4, 16'hD543,
 16'hAEB6, 16'hA451, 16'hA8A9, 16'hA55B,
 16'hA0A3, 16'hAB5E, 16'hB8A1, 16'hB35F,
 16'hA0A3, 16'h835A, 16'h8000, 16'h8053,
 16'h8000, 16'h804B, 16'h84BA, 16'h8940,
 16'h97C6, 16'hC336, 16'hF7CE, 16'h1D2E,
 16'h30D4, 16'h492B, 16'h5DD7, 16'h6F28,
 16'h79D8, 16'h7628, 16'h6BD7, 16'h582C,
 16'h3FD0, 16'h1F34, 16'hE4C8, 16'hA93C,
 16'h8000, 16'h8042, 16'h8000, 16'h8048,
 16'h8001, 16'h8048, 16'hB9B9, 16'hE744,
 16'h00C0, 16'h213B, 16'h3FCB, 16'h5A2F,
 16'h6ED8, 16'h721F, 16'h5CEC, 16'h3808,
 16'h2305, 16'h1CED, 16'h1D20, 16'h1ED4,
 16'h2338, 16'h20BD, 16'h014C, 16'hD0AD,
 16'hA558, 16'h90A5, 16'h875C, 16'h92A4,
 16'hA95B, 16'hBCA8, 16'hD952, 16'h0AB6,
 16'h323F, 16'h42CE, 16'h4D24, 16'h49EB,
 16'h3806, 16'h2109, 16'h18E7, 16'h1D29,
 16'h20C8, 16'h3546, 16'h3AAD, 16'h315F,
 16'h2396, 16'h1573, 16'h2085, 16'h4580,
 16'h757E, 16'h7F83, 16'h7E7E, 16'h7F7F,
 16'h7E85, 16'h7F74, 16'h7B96, 16'h625F,
 16'h2CAD, 16'hE947, 16'hA6C5, 16'h802E,
 16'h8000, 16'h8010, 16'h92FF, 16'hC6F4,
 16'hE517, 16'h04E0, 16'h2828, 16'h36D1,
 16'h2E35, 16'h22C6, 16'h0B3D, 16'hF0C3,
 16'hE33B, 16'hCCC9, 16'hAF31, 16'h9ED6,
 16'hA422, 16'hA8E9, 16'hA709, 16'hAB06,
 16'hCCEA, 16'hFD27, 16'h19C9, 16'h1546,
 16'hFFAA, 16'hDF67, 16'hC088, 16'hB988,
 16'hCE69, 16'hE3A4, 16'h0151, 16'h21B8,
 16'h2C40, 16'h40C7, 16'h5C34, 16'h76CF,
 16'h7E30, 16'h6BCF, 16'h3435, 16'hF3C4,
 16'hAF46, 16'h80AE, 16'h8001, 16'h8093,
 16'h927D, 16'hBA71, 16'hF2A2, 16'h2B4A,
 16'h57CA, 16'h5823, 16'h30EF, 16'hF700,
 16'hC310, 16'hAAE2, 16'hA72B, 16'h9EC9,
 16'h9842, 16'h90B5, 16'h8C51, 16'h8EAC,
 16'h9B54, 16'hCEB1, 16'h1546, 16'h61C5,
 16'h7F2D, 16'h7EE4, 16'h7F0A, 16'h7F0A,
 16'h7EDE, 16'h7F3D, 16'h7EA8, 16'h7073,
 16'h4E72, 16'h1DA8, 16'hCC3F, 16'h83D9,
 16'h8000, 16'h8105, 16'h8000, 16'h8126,
 16'h8000, 16'h813A, 16'hA7C1, 16'hC940,
 16'hCDC2, 16'hC439, 16'hC1D0, 16'hE024,
 16'hF1EB, 16'hFE02, 16'hFF13, 16'hF8D6,
 16'hFC43, 16'h13A2, 16'h3B7A, 16'h5E6A,
 16'h7EB1, 16'h7F35, 16'h7EE5, 16'h7F01,
 16'h7F18, 16'h7ED0, 16'h7946, 16'h7EA7,
 16'h7F69, 16'h7E8B, 16'h7F7E, 16'h7E7B,
 16'h4A8A, 16'h0B72, 16'hD591, 16'h9C6F,
 16'h8090, 16'h8000, 16'h8088, 16'h8001,
 16'h807D, 16'hAD89, 16'hF171, 16'h0094,
 16'hF167, 16'hCE9F, 16'hA95B, 16'h90AB,
 16'h9B50, 16'hBCB4, 16'hCF48, 16'hDBBC,
 16'hE741, 16'hE6C3, 16'hEA38, 16'hF2CC,
 16'hFD30, 16'h19D5, 16'h5425, 16'h7EE2,
 16'h7F16, 16'h7EF3, 16'h7F03, 16'h7F09,
 16'h7EE9, 16'h5E26, 16'h22CA, 16'hF347,
 16'hD4A8, 16'hE068, 16'hFF87, 16'h238B,
 16'h3F63, 16'h4FAE, 16'h4241, 16'h0FD0,
 16'hC721, 16'h80EC, 16'h8000, 16'h8104,
 16'h8000, 16'h8112, 16'h8000, 16'h8116,
 16'h8000, 16'hB60F, 16'h05F8, 16'h49FF,
 16'h7E0B, 16'h7FE9, 16'h7E25, 16'h7FCB,
 16'h7E47, 16'h5EA5, 16'h3670, 16'h1079,
 16'hE99D, 16'hBF4E, 16'h8000, 16'h8024,
 16'h8000, 16'h8003, 16'h801B, 16'h8000,
 16'h8042, 16'h9CAD, 16'h0562, 16'h3F91,
 16'h547B, 16'h4E7A, 16'h5890, 16'h7468,
 16'h7F9E, 16'h7E5E, 16'h7FA4, 16'h785C,
 16'h53A2, 16'h4C62, 16'h5D98, 16'h7970,
 16'h7F88, 16'h7E80, 16'h7F77, 16'h7E93,
 16'h5462, 16'h0BAB, 16'hEA47, 16'hE8C7,
 16'h072C, 16'h26E0, 16'h4315, 16'h59F6,
 16'h57FE, 16'h400E, 16'h23E7, 16'h0723,
 16'hF2D5, 16'hE930, 16'hDFCC, 16'hDC37,
 16'hDEC8, 16'hE737, 16'hECCB, 16'hF731,
 16'hF2D4, 16'hD525, 16'hAEE4, 16'h8F13,
 16'h8EF7, 16'hAEFE, 16'hD70D, 16'hF2E6,
 16'h072A, 16'h14C6, 16'h1F49, 16'h3BA9,
 16'h6863, 16'h7E92, 16'h7F78, 16'h7E7F,
 16'h7F8A, 16'h7E6E, 16'h7F98, 16'h7E63,
 16'h7FA2, 16'h7E5B, 16'h37A5, 16'hE95D,
 16'hB7A0, 16'h9065, 16'h9B94, 16'hB974,
 16'hD783, 16'h0087, 16'h2E6E, 16'h599E,
 16'h6F55, 16'h56B9, 16'h2139, 16'hDED5,
 16'h9F1D, 16'h8000, 16'h8003, 16'h800E,
 16'h81E5, 16'h9127, 16'hA6CF, 16'hD739,
 16'h00C2, 16'h1341, 16'h1CBD, 16'h2844,
 16'h36BC, 16'h3C43, 16'h27BF, 16'hF33D,
 16'hC0CA, 16'h9F2D, 16'h9CDD, 16'hA118,
 16'h9CF3, 16'hA402, 16'hB509, 16'hBCEC,
 16'hC11F, 16'hC5D7, 16'hD531, 16'hDBC7,
 16'hD240, 16'hD1BC, 16'hCB47, 16'hB9B6,
 16'hA94A, 16'hAFB8, 16'hBA46, 16'hC7BE,
 16'hE73C, 16'h14CB, 16'h402D, 16'h64DC,
 16'h6F19, 16'h61F4, 16'h48FF, 16'h240E,
 16'h0FE6, 16'h0F24, 16'h12D3, 16'h0937,
 16'hF6BF, 16'hE749, 16'hD6B0, 16'hD556,
 16'hF2A6, 16'h215E, 16'h5C9D, 16'h7F65,
 16'h7E9C, 16'h7662, 16'h6BA2, 16'h5A59,
 16'h4FAC, 16'h374E, 16'h15B9, 16'h003F,
 16'hEECA, 16'hE52E, 16'hDBD9, 16'hE320,
 16'hF3E6, 16'h0714, 16'h0FF2, 16'h1508,
 16'h1CFE, 16'h22FD, 16'h2408, 16'h23F3,
 16'h2711, 16'h1EEC, 16'h1A15, 16'h19EC,
 16'h2313, 16'h2CEE, 16'h3710, 16'h3AF3,
 16'h3B0A, 16'h3EF9, 16'h3B04, 16'h30FF,
 16'h26FE, 16'h2106, 16'h15F5, 16'h0910,
 16'hF6EB, 16'hEA1A, 16'hE4E2, 16'hE321,
 16'hE2DC, 16'hE026, 16'hE6D9, 16'hE928,
 16'hE2D7, 16'hDC29, 16'hCED9, 16'hC625,
 16'hC5DC, 16'hC722, 16'hCAE0, 16'hCD1E,
 16'hCCE7, 16'hD212, 16'hE4F4, 16'hFB06,
 16'h0900, 16'h0FFB, 16'h1A0A, 16'h22F1,
 16'h2E14, 16'h30E6, 16'h2D20, 16'h2CDA,
 16'h212D, 16'h18CC, 16'h0938, 16'hEEC6,
 16'hD23B, 16'hB4C5, 16'h9D3A, 16'h95C8,
 16'h9D36, 16'hA4CD, 16'hBA2F, 16'hD6D6,
 16'hEA25, 16'hF6E1, 16'h0517, 16'h14F1,
 16'h2308, 16'h2CFF, 16'h2DF9, 16'h2410,
 16'h12E5, 16'h0927, 16'h06CE, 16'h053B,
 16'h06BC, 16'h0B4D, 16'h06AB, 16'hF85C,
 16'hDE9E, 16'hC865, 16'hC09A, 16'hBA67,
 16'hC097, 16'hCB6A, 16'hD496, 16'hE369,
 16'hF69B, 16'h0260, 16'h0BA4, 16'h1357,
 16'h0EB0, 16'h0749, 16'h08BF, 16'h1938,
 16'h27D1, 16'h2826, 16'h2AE4, 16'h2111,
 16'h0AFA, 16'hFAFB, 16'hEA0F, 16'hF0E9,
 16'h071E, 16'h2ADB, 16'h4F2C, 16'h6ACD,
 16'h7F39, 16'h7EC2, 16'h7F41, 16'h7EBF,
 16'h7F41, 16'h5CBE, 16'h1A42, 16'hCCBF,
 16'h913F, 16'h8002, 16'h8338, 16'hADCC,
 16'hCF30, 16'hDAD4, 16'hE727, 16'hF7DF,
 16'h001A, 16'hF6ED, 16'hF10C, 16'hDBFB,
 16'hC5FE, 16'hB309, 16'h9EF0, 16'h9117,
 16'h86E1, 16'h8C27, 16'h9AD2, 16'hB034,
 16'hD0C8, 16'h023A, 16'h3AC4, 16'h543E,
 16'h49C0, 16'h2B42, 16'h0ABC, 16'hF145,
 16'hE9BC, 16'hF442, 16'hF6C1, 16'h013C,
 16'h0BC6, 16'h0C39, 16'h18C8, 16'h2B36,
 16'h3ECE, 16'h432E, 16'h2CD5, 16'h0227,
 16'hDBDD, 16'hB920, 16'h96E4, 16'h8D18,
 16'h95EB, 16'hA411, 16'hB9F4, 16'hE307,
 16'h0EFD, 16'h3100, 16'h3704, 16'h1CF6,
 16'hF711, 16'hD4E7, 16'hC722, 16'hCCD7,
 16'hD92F, 16'hDACA, 16'hCF3E, 16'hC6BA,
 16'hC74F, 16'hCEA6, 16'hF766, 16'h2A8D,
 16'h5881, 16'h7E70, 16'h7F9E, 16'h7855,
 16'h6CB8, 16'h603C, 16'h53CF, 16'h4926,
 16'h3FE5, 16'h2C10, 16'h0FFA, 16'hD0FE,
 16'h9409, 16'h8000, 16'h8114, 16'h8000,
 16'h8119, 16'h8000, 16'h8111, 16'hACF6,
 16'hC902, 16'hCE07, 16'hC3EE, 16'hC520,
 16'hDFD0, 16'hF042, 16'hFBAB, 16'hFA68,
 16'hF883, 16'hFA93, 16'h1057, 16'h31C0,
 16'h4D28, 16'h6FEF, 16'h7EFA, 16'h7F1C,
 16'h7ECF, 16'h7F45, 16'h75A8, 16'h6C6B,
 16'h7583, 16'h7F8C, 16'h7E67, 16'h7FA5,
 16'h7B51, 16'h4DB7, 16'h1543, 16'hE5C1,
 16'hAA3E, 16'h80C1, 16'h8002, 16'h80BD,
 16'h8002, 16'h80B4, 16'hAF52, 16'hEDA7,
 16'hFA60, 16'hE998, 16'hC671, 16'hA486,
 16'h8E83, 16'h9874, 16'hB995, 16'hCD61,
 16'hDEAB, 16'hE74A, 16'hE4BF, 16'hEA38,
 16'hF0D2, 16'h0024, 16'h19E8, 16'h540B,
 16'h7F00, 16'h7EF5, 16'h7F18, 16'h7EDB,
 16'h7F32, 16'h7EC0, 16'h5E4E, 16'h22A3,
 16'hF36D, 16'hD483, 16'hE08D, 16'hFF63,
 16'h23AD, 16'h3F43, 16'h4FCB, 16'h4228,
 16'h0FE5, 16'hC710, 16'h80F9, 16'h8000,
 16'h8106, 16'h8000, 16'h810D, 16'h8000,
 16'h810D, 16'h8000, 16'hB604, 16'h0604,
 16'h49F2, 16'h7E1A, 16'h7FDA, 16'h7E34,
 16'h7FBC, 16'h7E54, 16'h5E9B, 16'h3678,
 16'h1074, 16'hE9A1, 16'hBF49, 16'h8000,
 16'h801D, 16'h8000, 16'h8000, 16'h801E,
 16'h8000, 16'h8042, 16'h9CAF, 16'h055D,
 16'h3F98, 16'h5472, 16'h4E86, 16'h5881,
 16'h7478, 16'h7F8C, 16'h7E72, 16'h7F8F,
 16'h7873, 16'h5389, 16'h4C7A, 16'h5D82,
 16'h7983, 16'h7F78, 16'h7E8E, 16'h7F6B,
 16'h7E9D, 16'h545B, 16'h0BAD, 16'hEA4B,
 16'hE8BC, 16'h073E, 16'h26C8, 16'h4332,
 16'h59D5, 16'h5824, 16'h3FE2, 16'h2419,
 16'h06EB, 16'hF312, 16'hE8F0, 16'hE00E,
 16'hDBF4, 16'hDF0B, 16'hE6F5, 16'hED0B,
 16'hF6F5, 16'hF30B, 16'hD4F4, 16'hAB0E,
 16'h8CF0, 16'h8C12, 16'hADEC, 16'hD515,
 16'hF2EB, 16'h0516, 16'h14E8, 16'h211A,
 16'h3BE3, 16'h6C21, 16'h7EDB, 16'h7F29,
 16'h7ED3, 16'h7F30, 16'h7ECE, 16'h7F34,
 16'h7EC9, 16'h7F39, 16'h7EC6, 16'h3F3C,
 16'hE9C2, 16'hB33F, 16'h8CBF, 16'h9644,
 16'hB2BB, 16'hD245, 16'hFCBB, 16'h3144,
 16'h61BF, 16'h7A3E, 16'h60C5, 16'h2437,
 16'hDFCE, 16'h962C, 16'h8001, 16'h801F,
 16'h8002, 16'h8014, 16'h8000, 16'h980B,
 16'hCCFA, 16'hFD00, 16'h1006, 16'h1CF5,
 16'h270F, 16'h36EF, 16'h4011, 16'h27F0,
 16'hF10E, 16'hB4F5, 16'h9307, 16'h90FF,
 16'h97FA, 16'h930D, 16'h97EC, 16'hAF1B,
 16'hB8DE, 16'hB929, 16'hB8D0, 16'hC837,
 16'hD0C2, 16'hC844, 16'hC5B6, 16'hBA50,
 16'hA0AC, 16'h8C57, 16'h92A6, 16'hA55A,
 16'hB8A9, 16'hE353, 16'h1EB3, 16'h5846,
 16'h7EC1, 16'h7F37, 16'h78D2, 16'h5824,
 16'h2AE7, 16'h150D, 16'h12FF, 16'h12F5,
 16'h0517, 16'hE6DE, 16'hCD2D, 16'hB6C8,
 16'hB542, 16'hDBB5, 16'h1D54, 16'h6FA4,
 16'h7F64, 16'h7E95, 16'h7F70, 16'h7E8D,
 16'h7F75, 16'h7E8A, 16'h7A76, 16'h4F8A,
 16'h2D75, 16'h148D, 16'hFB70, 16'hE494,
 16'hE567, 16'hF29E, 16'h075D, 16'h12A7,
 16'h1656, 16'h18AD, 16'h1550, 16'h12B4,
 16'h1047, 16'h14BE, 16'h0C3E, 16'h0EC4,
 16'h0F3D, 16'h0FC1, 16'h0C3F, 16'h0BC2,
 16'h103D, 16'h0BC4, 16'h0F3C, 16'h0EC1,
 16'h0F44, 16'h0EB8, 16'h0B4B, 16'h0BB3,
 16'h0C4E, 16'h0BB1, 16'h0C52, 16'h08AA,
 16'h075A, 16'h08A2, 16'h0962, 16'h089B,
 16'h0568, 16'h0195, 16'h016C, 16'h0196,
 16'h0166, 16'h009E, 16'h005F, 16'hFFA4,
 16'hFD59, 16'hFCAB, 16'hFD4E, 16'hFFBB,
 16'h003D, 16'hFFCB, 16'hF82C, 16'hF7DE,
 16'hF718, 16'hFAF2, 16'hF705, 16'hF402,
 16'hF7F7, 16'hF410, 16'hF6EA, 16'hF71C,
 16'hF6DF, 16'hF323, 16'hF6DB, 16'hF427,
 16'hF0D9, 16'hF327, 16'hF2D9, 16'hF324,
 16'hF2E1, 16'hF11A, 16'hECEB, 16'hEA10,
 16'hECF6, 16'hF104, 16'hED03, 16'hECF5,
 16'hED12, 16'hECE9, 16'hED1B, 16'hECE3,
 16'hED1E, 16'hECE0, 16'hED21, 16'hECDF,
 16'hF120, 16'hF0E3, 16'hEF18, 16'hF2EE,
 16'hF40B, 16'hF3FD, 16'hF2FB, 16'hF30E,
 16'hF0E8, 16'hE022, 16'hCCD5, 16'hCB32,
 16'hCACA, 16'hC339, 16'hC6C5, 16'hE93B,
 16'h18C7, 16'h3736, 16'h34CF, 16'h1A2C,
 16'hF7D8, 16'hD723, 16'hBCE5, 16'hB011,
 16'hADFB, 16'hAFF7, 16'hBF16, 16'hD6E0,
 16'h0F28, 16'h53D0, 16'h7F37, 16'h7EC4,
 16'h7F3F, 16'h7EC1, 16'h7F3B, 16'h6ACB,
 16'h0F2D, 16'hCCDE, 16'hBA13, 16'hC300,
 16'hDBEA, 16'hDC2F, 16'hCAB6, 16'hB966,
 16'hA47C, 16'h98A5, 16'h9039, 16'h8FE9,
 16'h87F5, 16'h812C, 16'h8000, 16'h8166,
 16'h8000, 16'h8198, 16'h8000, 16'h84BD,
 16'hC537, 16'h20D0, 16'h782E, 16'h7FFF,
 16'h7D37, 16'h7FFE, 16'h7D53, 16'h719A,
 16'h667B, 16'h666D, 16'h51AE, 16'h2C35,
 16'hFEEB, 16'hDFF2, 16'hC530, 16'hB7AF,
 16'hAD73, 16'hAB6D, 16'hA0B1, 16'h8331,
 16'h8002, 16'hA0FE, 16'hD117, 16'hF0D7,
 16'hEF39, 16'hDFB8, 16'hCD55, 16'hBCA1,
 16'hB567, 16'hB493, 16'hB971, 16'hCA8D,
 16'hE074, 16'hF78C, 16'h1573, 16'h308E,
 16'h5472, 16'h7E8C, 16'h7F76, 16'h7E88,
 16'h7F7B, 16'h7E81, 16'h7F84, 16'h7E75,
 16'h7F93, 16'h3665, 16'hEAA3, 16'hAA56,
 16'h80B2, 16'h8000, 16'h80C2, 16'h8000,
 16'h80CD, 16'h8000, 16'h85D2, 16'hC22D,
 16'hE3D2, 16'hE832, 16'hE7C7, 16'hDF41,
 16'hD9B5, 16'hD157, 16'hCD9D, 16'hCE70,
 16'hCD82, 16'hCE8A, 16'hD26C, 16'hD89F,
 16'hDC56, 16'hE2B4, 16'hE742, 16'hECC7,
 16'hEF33, 16'hF2CF, 16'hF332, 16'hF3C9,
 16'hE540, 16'hB6B4, 16'h985A, 16'h8696,
 16'h877C, 16'h9770, 16'hB0A6, 16'hCA42,
 16'hF1D8, 16'h120E, 16'h2C0B, 16'h48DD,
 16'h5B3A, 16'h6AB0, 16'h7363, 16'h7D8E,
 16'h7FFF, 16'h7D7C, 16'h7FFF, 16'h7D7C,
 16'h7FFF, 16'h7D8D, 16'h7FFF, 16'h78B3,
 16'hEE34, 16'h87EA, 16'h80F5, 16'h8000,
 16'h80A9, 16'h8000, 16'h8054, 16'h96D9,
 16'hDFFA, 16'h0232, 16'hF7A4, 16'hD984,
 16'hB457, 16'h93CB, 16'h8216, 16'h8106,
 16'h8003, 16'h8131, 16'h8003, 16'h844B,
 16'h8DAF, 16'h9953, 16'h96AE, 16'h814B,
 16'h8000, 16'h8A32, 16'hBBE1, 16'hEE09,
 16'hFC0E, 16'hF8DA, 16'hE83F, 16'hE5A8,
 16'h0171, 16'h3277, 16'h61A0, 16'h754A,
 16'h64CC, 16'h461F, 16'h23F3, 16'h0AFE,
 16'hF40E, 16'hE6E9, 16'hE31F, 16'hDBDB,
 16'hDF28, 16'hE2D7, 16'hE027, 16'hD8DF,
 16'hBD1A, 16'hA3EE, 16'h9607, 16'h9F04,
 16'hD6F1, 16'h1F1C, 16'h4ED7, 16'h5734,
 16'h49C0, 16'h2E4C, 16'h27A9, 16'h3161,
 16'h2A96, 16'h1A72, 16'h0488, 16'h017D,
 16'h157D, 16'h1A88, 16'h1976, 16'h1D8B,
 16'h3676, 16'h5A86, 16'h647E, 16'h617F,
 16'h5C85, 16'h6175, 16'h5692, 16'h3266,
 16'h04A4, 16'hD952, 16'hB8B7, 16'h9D3F,
 16'h8ECC, 16'h892A, 16'h8BE1, 16'h9114,
 16'h97F5, 16'h9F02, 16'hA908, 16'hAAEF,
 16'h9D19, 16'hA4DF, 16'hB327, 16'hBED5,
 16'hDC2F, 16'h04CC, 16'h1A38, 16'h14C5,
 16'h133D, 16'h06C4, 16'hFD38, 16'hFACD,
 16'hF32D, 16'hF0DA, 16'hEF1E, 16'hECEB,
 16'hE90B, 16'hE9FF, 16'hE8F7, 16'hD913,
 16'hD6E2, 16'hF32B, 16'h08C7, 16'h1546,
 16'h14AE, 16'h105C, 16'h0E9C, 16'h096B,
 16'h048E, 16'h0179, 16'hFF81, 16'hFD83,
 16'hFC7C, 16'hFB83, 16'hFF80, 16'hFD7B,
 16'hFF8B, 16'h006E, 16'hFF9A, 16'h005E,
 16'h01AA, 16'h004D, 16'hFFBC, 16'hFD3B,
 16'hFCCE, 16'h012A, 16'h00DD, 16'h021B,
 16'h04EE, 16'h010A, 16'hFFFD, 16'hFFFD,
 16'hFD07, 16'hFCF7, 16'hF109, 16'hF0F9,
 16'hED04, 16'hF300, 16'h04FB, 16'h0F08,
 16'h14F5, 16'h100F, 16'h08ED, 16'h0717,
 16'h00E4, 16'hF820, 16'hFADD, 16'hF125,
 16'hE9DB, 16'hF124, 16'hF6DD, 16'hF722,
 16'hFAE0, 16'hF81C, 16'hF7EA, 16'hF70F,
 16'hF2F8, 16'hF702, 16'hF402, 16'hF0FB,
 16'hE709, 16'hCAF2, 16'hBA13, 16'hC7E9,
 16'hF11A, 16'h14E5, 16'h241B, 16'h36E6,
 16'h3C18, 16'h34EB, 16'h2310, 16'h0EF8,
 16'hFFFF, 16'hF409, 16'hEEEF, 16'hE71A,
 16'hE6DD, 16'hE72C, 16'hE2C9, 16'hE743,
 16'hE8B3, 16'hE956, 16'hE9A1, 16'hEA66,
 16'hEC95, 16'hED6F, 16'hF08F, 16'hEF72,
 16'hF28D, 16'hF473, 16'hF38F, 16'hF46E,
 16'hF697, 16'hF463, 16'hF7A3, 16'hF758,
 16'hF6AE, 16'hF74B, 16'hF6BD, 16'hF73B,
 16'hF6CC, 16'hF12F, 16'hD4D4, 16'hB72A,
 16'h9CD9, 16'hA124, 16'hC5DD, 16'hE723,
 16'hFCDC, 16'h0726, 16'h0BD7, 16'h092C,
 16'h06D1, 16'h0733, 16'h0BC8, 16'h2B3C,
 16'h4FBF, 16'h6C47, 16'h7EB3, 16'h7F53,
 16'h7EA8, 16'h7F5A, 16'h71A6, 16'h4A5A,
 16'h2AA8, 16'h0154, 16'hD6B1, 16'hC749,
 16'hC2BE, 16'hB73B, 16'hA8CD, 16'hB029,
 16'hCCE3, 16'hF10F, 16'hF7FF, 16'hFCF3,
 16'h0B1B, 16'h0FD7, 16'h0736, 16'hE6BC,
 16'hC753, 16'hAA9F, 16'h986D, 16'h8E88,
 16'h8582, 16'h8000, 16'h8091, 16'h8000,
 16'h8096, 16'h926B, 16'hA592, 16'hC272,
 16'hF18A, 16'h2D7C, 16'h627C, 16'h748D,
 16'h6568, 16'h52A6, 16'h314A, 16'h14C7,
 16'h0128, 16'hEEEA, 16'hEA04, 16'hDF0D,
 16'hDFE2, 16'hE32E, 16'hE6C3, 16'hED4C,
 16'hF2A6, 16'hF767, 16'hF78C, 16'hE380,
 16'hC675, 16'hCD94, 16'hD866, 16'hDF9D,
 16'hE462, 16'hE99E, 16'h0863, 16'h3B9B,
 16'h6F68, 16'h7F93, 16'h7475, 16'h5381,
 16'h378A, 16'h326B, 16'h2DA0, 16'h2355,
 16'h18B5, 16'h2340, 16'h44CD, 16'h5A27,
 16'h57E4, 16'h5811, 16'h60F9, 16'h60FD,
 16'h4A0E, 16'h1EE8, 16'hF821, 16'hDED7,
 16'hBF2F, 16'hAFCC, 16'hAB39, 16'hA6C2,
 16'hAB42, 16'hAFBC, 16'hB545, 16'hBCBB,
 16'hC344, 16'hC6BD, 16'hCF42, 16'hD4BF,
 16'hD940, 16'hDAC2, 16'hDC3B, 16'hD6C8,
 16'hBD34, 16'hA3D0, 16'h932C, 16'h8BD8,
 16'h9323, 16'hA0E2, 16'hC71A, 16'h00EA,
 16'h2811, 16'h3FF3, 16'h4609, 16'h4CFD,
 16'h67FD, 16'h7F07, 16'h7EF5, 16'h7F0F,
 16'h7EED, 16'h7F18, 16'h7EE2, 16'h5E23,
 16'h3FD9, 16'h2B2C, 16'h0BCF, 16'hDC36,
 16'hAEC4, 16'h9142, 16'h8000, 16'h8049,
 16'h8000, 16'h804F, 16'h8000, 16'h8054,
 16'h96AA, 16'hBF57, 16'hE2A9, 16'hEF56,
 16'hECAB, 16'hDC54, 16'hCAAE, 16'hCB4E,
 16'hE6B7, 16'h1A43, 16'h3FC5, 16'h4A32,
 16'h3BD8, 16'h321D, 16'h2AEF, 16'h1A05,
 16'h2306, 16'h31EF, 16'h461C, 16'h52D9,
 16'h3833, 16'h0AC0, 16'hD14C, 16'h9AA9,
 16'h8F62, 16'h8B94, 16'h9375, 16'hB483,
 16'hE083, 16'h0E7A, 16'h1F87, 16'h197A,
 16'h0583, 16'hF282, 16'hDC78, 16'hC290,
 16'hB365, 16'hADA7, 16'hA14D, 16'h96C1,
 16'h8C31, 16'h8CDC, 16'h9716, 16'hA6F8,
 16'hDAFB, 16'h2311, 16'h61E4, 16'h7F27,
 16'h7ECE, 16'h7F3C, 16'h7EBB, 16'h7F4B,
 16'h7EB2, 16'h7250, 16'h4CB0, 16'h1A4F,
 16'hFCB2, 16'hE74B, 16'hDEBA, 16'hE041,
 16'hFAC5, 16'h1635, 16'h20D1, 16'h132A,
 16'hFCDA, 16'hED21, 16'hDAE5, 16'hD516,
 16'hCEEF, 16'hCF0D, 16'hCEF5, 16'hD50A,
 16'hD4F7, 16'hDB09, 16'hDFF6, 16'hE50B,
 16'hE8F2, 16'hED13, 16'hF0E9, 16'hF31A,
 16'hFAE3, 16'hF820, 16'hFADC, 16'h0029,
 16'h01D2, 16'hF733, 16'hDFC8, 16'hBA3D,
 16'hA3BD, 16'h934A, 16'h96AF, 16'hA757,
 16'hBEA3, 16'hD963, 16'hF698, 16'h166D,
 16'h2D8D, 16'h467A, 16'h5D7F, 16'h7F89,
 16'h7E6D, 16'h7F9D, 16'h7E59, 16'h7FB2,
 16'h7E43, 16'h7FC7, 16'h782E, 16'h28DD,
 16'hFF19, 16'hEFF0, 16'hDE07, 16'hE602,
 16'hF9F7, 16'h170E, 16'h26ED, 16'h1B18,
 16'hFEE4, 16'hE01F, 16'hAEE0, 16'h831F,
 16'h8003, 16'h8119, 16'h8002, 16'h810F,
 16'h8001, 16'h8DFF, 16'hB80A, 16'hDCEC,
 16'h0120, 16'h16D4, 16'h1438, 16'h09BC,
 16'h014F, 16'h07A6, 16'hF767, 16'hDC8C,
 16'hC781, 16'hB572, 16'hA899, 16'hA15D,
 16'hA3AD, 16'hA14A, 16'h95BD, 16'h913C,
 16'hAFCB, 16'hDB2E, 16'h00D9, 16'h1020,
 16'h0FE7, 16'h1512, 16'h12F4, 16'h1306,
 16'h0F01, 16'h0BF9, 16'h0C0C, 16'h0AEE,
 16'h0C18, 16'h0EE2, 16'h1525, 16'h14D4,
 16'h1632, 16'h18C9, 16'h1A3A, 16'h1CC4,
 16'h1D3E, 16'h1EBF, 16'h2145, 16'h20B7,
 16'h214D, 16'h20B0, 16'h2150, 16'h20B2,
 16'h1D4C, 16'h20B7, 16'h1D46, 16'h18BC,
 16'h1941, 16'h15C4, 16'h1536, 16'h12D1,
 16'h1027, 16'h12E2, 16'h0C15, 16'h06F4,
 16'hF302, 16'hCF08, 16'hB4EE, 16'h9F1C,
 16'h9ADB, 16'hA52E, 16'hB6C9, 16'hCD3F,
 16'hE8B9, 16'h054F, 16'h30AA, 16'h685D,
 16'h7E9D, 16'h7F67, 16'h7E96, 16'h7F6C,
 16'h7E93, 16'h7F6E, 16'h7E92, 16'h546B,
 16'h199A, 16'hE560, 16'hC0A6, 16'hB954,
 16'hD0B2, 16'h0047, 16'h2DC2, 16'h5734,
 16'h6AD6, 16'h671F, 16'h44ED, 16'h0107,
 16'hBA05, 16'h8CEF, 16'h801D, 16'h8000,
 16'h8035, 16'h8000, 16'h8049, 16'h8000,
 16'h805A, 16'h8000, 16'hB367, 16'h0693,
 16'h4671, 16'h788D, 16'h7C74, 16'h648E,
 16'h4D6D, 16'h3B99, 16'h235F, 16'hFFAB,
 16'hE04B, 16'hC5C0, 16'hB534, 16'hADD9,
 16'hAB18, 16'hADFA, 16'hB4F3, 16'hBD21,
 16'hB8CA, 16'hB34A, 16'hB8A3, 16'hB56F,
 16'hB281, 16'hB58E, 16'hB863, 16'hCFAC,
 16'hFC45, 16'h35C9, 16'h5C2C, 16'h65DD,
 16'h601C, 16'h53E8, 16'h5216, 16'h62EB,
 16'h7E18, 16'h7FE2, 16'h7E25, 16'h7FD1,
 16'h753B, 16'h50BA, 16'h2352, 16'h02A0,
 16'hF36E, 16'hFD82, 16'h0490, 16'h055F,
 16'h08B2, 16'h163C, 16'h27D6, 16'h2817,
 16'h18FB, 16'h06F6, 16'hF318, 16'hE8DB,
 16'hDC31, 16'hD6C2, 16'hD94B, 16'hD8AA,
 16'hDF5F, 16'hE49A, 16'hE76C, 16'hEC8F,
 16'hF175, 16'hF388, 16'hF379, 16'hF388,
 16'hFD76, 16'h048D, 16'h056E, 16'hFF99,
 16'hF35F, 16'hE6AA, 16'hEF4C, 16'hFFBF,
 16'h0B35, 16'h14D8, 16'h161A, 16'h15F5,
 16'h0FFC, 16'h1014, 16'h0ADB, 16'h0F35,
 16'h18BC, 16'h2352, 16'h2DA2, 16'h3869,
 16'h488B, 16'h4A81, 16'h4274, 16'h3296,
 16'h2261, 16'h16A7, 16'h0A52, 16'hF8B4,
 16'hF348, 16'hF1B9, 16'hEC48, 16'hE5B6,
 16'hE64C, 16'hF1B2, 16'h0051, 16'h05A9,
 16'h045F, 16'h0999, 16'h0A6F, 16'h0288,
 16'hF681, 16'hEA77, 16'hDB92, 16'hD266,
 16'hC0A0, 16'hA959, 16'hA6AF, 16'hAB4A,
 16'hB8BD, 16'hC63D, 16'hC0C8, 16'hC133,
 16'hD1D1, 16'hEF2C, 16'h0BD7, 16'h2827,
 16'h2CDB, 16'h2322, 16'h20E2, 16'h1F19,
 16'h34EB, 16'h3C12, 16'h3BF1, 16'h3F0C,
 16'h3FF6, 16'h3B07, 16'h23FD, 16'h08FF,
 16'hEA04, 16'hDAF8, 16'hD70E, 16'hD6EC,
 16'hD118, 16'hD1E5, 16'hE71E, 16'hEEDF,
 16'hE524, 16'hDFD9, 16'hDF2A, 16'hE6D3,
 16'hFB2E, 16'h0AD3, 16'h0C2B, 16'h01D9,
 16'hF322, 16'hE4E2, 16'hEA1A, 16'hF3EC,
 16'h000D, 16'h19FC, 16'h42F9, 16'h7012,
 16'h7EE3, 16'h7F29, 16'h78CA, 16'h7244,
 16'h6AAD, 16'h5363, 16'h238C, 16'hF784,
 16'hDB6D, 16'hC1A2, 16'hAA50, 16'h91BE,
 16'h8833, 16'h85DB, 16'h8819, 16'h89F1,
 16'h9508, 16'hA9FD, 16'hC4FE, 16'hE105,
 16'hF2FA, 16'hF407, 16'hE7FA, 16'hE002,
 16'hD003, 16'hC7F5, 16'hC616, 16'hC1DE,
 16'hBE2F, 16'hC8C2, 16'hD44E, 16'hE9A0,
 16'h0F74, 16'h2477, 16'h3A9E, 16'h464B,
 16'h4FCE, 16'h6719, 16'h7C00, 16'h7BE8,
 16'h6F2E, 16'h6ABC, 16'h6C5A, 16'h5D91,
 16'h4383, 16'h346B, 16'h28A4, 16'h184E,
 16'hF4BF, 16'hD136, 16'hB9D3, 16'hA826,
 16'h9BDE, 16'h8C21, 16'h80DE, 16'h8824,
 16'h9DD8, 16'hB62E, 16'hD2CA, 16'hEE41,
 16'hF7B2, 16'hF65C, 16'hEA95, 16'hDE79,
 16'hDF7A, 16'hF394, 16'h195E, 16'h36B0,
 16'h3F41, 16'h31CD, 16'h2B27, 16'h27E4,
 16'h1A11, 16'h1EFA, 16'h2DFC, 16'h3C0C,
 16'h42EF, 16'h3114, 16'h0EEB, 16'hDC14,
 16'hB2ED, 16'hA912, 16'hA4F1, 16'hA90A,
 16'hBEFD, 16'hDFFA, 16'h0210, 16'h14E5,
 16'h1025, 16'h06D2, 16'h0038, 16'hF0BC,
 16'hDB51, 16'hCEA2, 16'hC66A, 16'hB88C,
 16'hAE7A, 16'hA083, 16'h9F80, 16'hAA7E,
 16'hBA83, 16'hE87D, 16'h2482, 16'h5681,
 16'h757A, 16'h7E8D, 16'h7F6B, 16'h749F,
 16'h6B55, 16'h6BB8, 16'h5D3A, 16'h3BD4,
 16'h101E, 16'hF6F1, 16'hE700, 16'hDB0E,
 16'hDFE4, 16'hFB28, 16'h12CF, 16'h1A3A,
 16'h0EBE, 16'hFB49, 16'hEEB0, 16'hDC56,
 16'hD6A7, 16'hD15A, 16'hD0A7, 16'hD157,
 16'hD4AB, 16'hD753, 16'hDBB1, 16'hE34A,
 16'hE6BB, 16'hEA3E, 16'hEECA, 16'hF12F,
 16'hF3D9, 16'hF81E, 16'hF7EA, 16'hFB0E,
 16'hFFFB, 16'hFFFB, 16'hF70F, 16'hE2E8,
 16'hBD21, 16'hA6D6, 16'h9731, 16'h9AC9,
 16'hA93D, 16'hBEBE, 16'hDB48, 16'hF6B0,
 16'h1559, 16'h2D9D, 16'h456E, 16'h5D87,
 16'h7F85, 16'h7E6F, 16'h7F9C, 16'h7E59,
 16'h7FB3, 16'h7E41, 16'h7FCB, 16'h7829,
 16'h28E3, 16'hFF12, 16'hEFF8, 16'hDDFE,
 16'hE60B, 16'hF9EE, 16'h1718, 16'h26E2,
 16'h1B22, 16'hFEDC, 16'hE026, 16'hAED9,
 16'h8325, 16'h8001, 16'h811C, 16'h8003,
 16'h810E, 16'h8003, 16'h8DFC, 16'hB80E,
 16'hDCE7, 16'h0125, 16'h16CF, 16'h143D,
 16'h09B8, 16'h0152, 16'h07A4, 16'hF766,
 16'hDC8F, 16'hC77E, 16'hB575, 16'hA897,
 16'hA15D, 16'hA3AE, 16'hA149, 16'h95BF,
 16'h913A, 16'hAFCD, 16'hDB2B, 16'h00DD,
 16'h101C, 16'h0FEB, 16'h150F, 16'h12F6,
 16'h1304, 16'h0F02, 16'h0BF9, 16'h0C0C,
 16'h0AEF, 16'h0C16, 16'h0EE5, 16'h151F,
 16'h14DD, 16'h1628, 16'h18D3, 16'h1A33,
 16'h1CC7, 16'h1D3D, 16'h1EC1, 16'h2140,
 16'h20BF, 16'h2143, 16'h20BB, 16'h2147,
 16'h20B9, 16'h1D45, 16'h20BD, 16'h1D41,
 16'h18C2, 16'h193B, 16'h15C9, 16'h1531,
 16'h12D6, 16'h1024, 16'h12E1, 16'h0C19,
 16'h06EE, 16'hF30B, 16'hCEFE, 16'hB4F8,
 16'h9F11, 16'h9AE6, 16'hA124, 16'hB4D2,
 16'hCB38, 16'hE6BE, 16'h074B, 16'h30AD,
 16'h685B, 16'h7E9D, 16'h7F6B, 16'h7E8D,
 16'h7F7B, 16'h7E7F, 16'h7F85, 16'h7E79,
 16'h5787, 16'h1C7A, 16'hE385, 16'hBC7D,
 16'hB780, 16'hCE84, 16'h0176, 16'h3192,
 16'h5A64, 16'h6FA7, 16'h6F4D, 16'h48C0,
 16'hFD32, 16'hB4DD, 16'h8214, 16'h8000,
 16'h8000, 16'h8019, 16'h8001, 16'h8033,
 16'h8001, 16'h8048, 16'h8000, 16'hA758,
 16'h08A4, 16'h535E, 16'h7EA3, 16'h7F59,
 16'h6FAD, 16'h544B, 16'h3FBF, 16'h2436,
 16'hFCD7, 16'hDF19, 16'hB9F8, 16'hA8F6,
 16'h9F1E, 16'h9CCE, 16'hA146, 16'hA8A6,
 16'hB36D, 16'hAA81, 16'hA790, 16'hAD60,
 16'hA5B0, 16'hA442, 16'hA7C8, 16'hAA31,
 16'hC6D3, 16'hFC2C, 16'h43D4, 16'h792E,
 16'h7FCD, 16'h7E3B, 16'h6BBB, 16'h6150,
 16'h70A3, 16'h7E6C, 16'h7F85, 16'h7E8B,
 16'h7F64, 16'h7EAC, 16'h6843, 16'h30CF,
 16'h0720, 16'hF7F0, 16'h0201, 16'h0C0B,
 16'h0BEB, 16'h151D, 16'h23DD, 16'h3C27,
 16'h3ED6, 16'h272C, 16'h0ED4, 16'hF42A,
 16'hE2DA, 16'hD220, 16'hCEE7, 16'hCF11,
 16'hCCF8, 16'hD4FF, 16'hDB0A, 16'hDFED,
 16'hE71B, 16'hEEDD, 16'hF12B, 16'hF0CE,
 16'hF338, 16'hFFC3, 16'h0B41, 16'h0EBB,
 16'h1049, 16'h0BB4, 16'h054E, 16'h0FB2,
 16'h164D, 16'h1CB5, 16'h1F48, 16'h1EBA,
 16'h1A44, 16'h14C0, 16'h133D, 16'h0BC5,
 16'h0F38, 16'h0BCA, 16'h0B35, 16'h0BCC,
 16'h0934, 16'h0ACB, 16'h0B35, 16'h0BCC,
 16'h0C34, 16'h08CB, 16'h0B36, 16'h0BC9,
 16'h0B38, 16'h0BC8, 16'h0C37, 16'h0ACA,
 16'h0735, 16'h0ACC, 16'h0732, 16'h08D0,
 16'h092D, 16'h08D7, 16'h0525, 16'h01E0,
 16'h011B, 16'hFFE9, 16'h0112, 16'hFFF4,
 16'hFD08, 16'hE2FD, 16'hC5FD, 16'hCF07,
 16'hE6F6, 16'hF70E, 16'hF6EF, 16'hE313,
 16'hD6EA, 16'hDB18, 16'hECE8, 16'hF419,
 16'hF6E6, 16'hF11A, 16'hE9E5, 16'hF11C,
 16'h0FE5, 16'h4A1A, 16'h6FE8, 16'h7F16,
 16'h7EEB, 16'h7F15, 16'h7EEB, 16'h6116,
 16'h27E9, 16'hE917, 16'hC0E9, 16'hB918,
 16'hB4E6, 16'hBA1D, 16'hDBDF, 16'hFD25,
 16'h04D7, 16'hEA2D, 16'hD4CF, 16'hCF34,
 16'hC2CA, 16'hB037, 16'h96C9, 16'h8736,
 16'h8002, 16'h8034, 16'h86CF, 16'h962C,
 16'hAADC, 16'hD21A, 16'h19F1, 16'h6103,
 16'h7F0A, 16'h7EE9, 16'h7F25, 16'h7ECC,
 16'h7F45, 16'h75A9, 16'h5D69, 16'h2786,
 16'hF78B, 16'hDE64, 16'hC3AD, 16'h9C42,
 16'h80CE, 16'h8000, 16'h80E8, 16'h8000,
 16'h80FD, 16'h8000, 16'h810A, 16'hBBF2,
 16'hFE11, 16'h21EC, 16'h1B15, 16'hFEED,
 16'hDC0F, 16'hC6F7, 16'hDA01, 16'hFC08,
 16'h10F0, 16'h1C17, 16'h2DE2, 16'h2725,
 16'h2BD4, 16'h2C35, 16'h1FC1, 16'h2749,
 16'h3FAD, 16'h575E, 16'h6598, 16'h5671,
 16'h2885, 16'h0685, 16'hFD72, 16'h0897,
 16'h095F, 16'h04AB, 16'h104B, 16'h23BF,
 16'h2B37, 16'h27D3, 16'h1F23, 16'h15E7,
 16'h0C0E, 16'h01FD, 16'hFFF9, 16'h0000,
 16'h11E5, 16'h0224, 16'h01D4, 16'h0733,
 16'h0BC6, 16'h0B41, 16'h0FB9, 16'h0F4D,
 16'h0FAD, 16'h1558, 16'h15A3, 16'h1962,
 16'h199A, 16'h1569, 16'h1895, 16'h156C,
 16'h1494, 16'h156A, 16'h1498, 16'h1367,
 16'h129B, 16'h1063, 16'h0E9F, 16'h0F5E,
 16'h0BA6, 16'h0B56, 16'h04AF, 16'h004B,
 16'hFABC, 16'hE93D, 16'hD1C9, 16'hD231,
 16'hDFD5, 16'hEA24, 16'h06E5, 16'h2D11,
 16'h44F9, 16'h48FD, 16'h490D, 16'h37EA,
 16'h281F, 16'h1ED7, 16'h0B34, 16'h01C1,
 16'h0C4A, 16'h23AB, 16'h325E, 16'h2D9B,
 16'h196C, 16'h008D, 16'hED79, 16'hDA81,
 16'hCF85, 16'hC577, 16'hC18B, 16'hC275,
 16'hBF89, 16'hC27A, 16'hC182, 16'hC083,
 16'hCB77, 16'hDE90, 16'hE369, 16'hE89E,
 16'hE95B, 16'hE8AC, 16'hE94C, 16'hE6BE,
 16'hE738, 16'hE8D1, 16'hEA26, 16'hE4E3,
 16'hE915, 16'hE9F3, 16'hEA05, 16'hED00,
 16'hEEFD, 16'hED05, 16'hECFB, 16'hF104,
 16'hF2FD, 16'hF101, 16'hF403, 16'hF6F7,
 16'hF411, 16'hF7E6, 16'hF423, 16'hF6D5,
 16'hF832, 16'hF7C6, 16'hF843, 16'hF7B4,
 16'hF856, 16'hF7A0, 16'hFB68, 16'h0091,
 16'h0076, 16'hEC85, 16'hE57F, 16'hF07D,
 16'h0085, 16'hFF7B, 16'hE984, 16'hCE7F,
 16'hB37C, 16'hA88A, 16'hB76D, 16'hE69E,
 16'h1A57, 16'h36B5, 16'h383E, 16'h37CF,
 16'h4324, 16'h57E9, 16'h5A0A, 16'h4503,
 16'h22F0, 16'hF81D, 16'hD6D7, 16'hBF33,
 16'hB2C4, 16'hB344, 16'hB9B5, 16'hD551,
 16'h0BAB, 16'h5057, 16'h7EAA, 16'h7F53,
 16'h7EB1, 16'h7F49, 16'h7EBF, 16'h623A,
 16'h23CD, 16'hDF2A, 16'hAEE0, 16'h9816,
 16'h84F5, 16'h8000, 16'h800C, 16'h97EB,
 16'hC31D, 16'hDBDB, 16'hEA2C, 16'h00CF,
 16'h1535, 16'h0EC8, 16'h0039, 16'hF0C7,
 16'hD73A, 16'hCAC6, 16'hD137, 16'hE6CE,
 16'hF82B, 16'hFCDD, 16'hEF1B, 16'hDAEC,
 16'hC80E, 16'hB9F8, 16'hB301, 16'hB007,
 16'hAEF0, 16'hA71A, 16'hA4DC, 16'h9B2D,
 16'h8CCB, 16'h873D, 16'h88BB, 16'h934D,
 16'hAAAA, 16'hC15E, 16'hF39C, 16'h2D6A,
 16'h5D90, 16'h7A76, 16'h7E83, 16'h7F85,
 16'h7973, 16'h7F94, 16'h7E66, 16'h7FA0,
 16'h7E5A, 16'h7FAC, 16'h7E4E, 16'h7FB7,
 16'h7E44, 16'h7FC1, 16'h7E3B, 16'h40C8,
 16'h0636, 16'hCBCA, 16'h8C38, 16'h80C5,
 16'h8004, 16'h89BB, 16'hBE4B, 16'hF3AF,
 16'h2059, 16'h389D, 16'h316E, 16'h1386,
 16'hEE87, 16'hD26C, 16'hB8A2, 16'h9F4F,
 16'h8CC1, 16'h802F, 16'h8001, 16'h8013,
 16'h8000, 16'h8000, 16'h8013, 16'h8000,
 16'h8027, 16'hA0D1, 16'hBD37, 16'hCEC2,
 16'hDF43, 16'hE8BA, 16'hFD46, 16'h20BD,
 16'h433F, 16'h66C6, 16'h7F34, 16'h7ED3,
 16'h7A25, 16'h60E4, 16'h4013, 16'h23F6,
 16'h0F00, 16'h010B, 16'h06E9, 16'h2B23,
 16'h61D2, 16'h7F38, 16'h7EBF, 16'h7F49,
 16'h7EAF, 16'h7959, 16'h3FA1, 16'hFB63,
 16'hBE9A, 16'h8967, 16'h8005, 16'h8067,
 16'h8003, 16'h8063, 16'hA6A1, 16'hF159,
 16'h36B0, 16'h6C45, 16'h7EC7, 16'h7F2C,
 16'h6AE2, 16'h3110, 16'h01FE, 16'hDFF4,
 16'hCD1A, 16'hAED8, 16'h8336, 16'h8000,
 16'h804E, 16'h8000, 16'h8060, 16'h8000,
 16'h8067, 16'h8000, 16'hBD65, 16'h189F,
 16'h4D5A, 16'h53B0, 16'h4042, 16'h36CF,
 16'h431E, 16'h56F7, 16'h6BF2, 16'h7C26,
 16'h6AC1, 16'h4959, 16'h2C8D, 16'h1D8C,
 16'h065C, 16'hDBBB, 16'hB431, 16'hA7E0,
 16'hA411, 16'h9FFC, 16'h99FA, 16'h990D,
 16'h9BF0, 16'hB80F, 16'hEDF6, 16'h3800,
 16'h7E0E, 16'h7FE1, 16'h7E35, 16'h7FB2,
 16'h7E69, 16'h7679, 16'h75A7, 16'h6838,
 16'h44EA, 16'h15F5, 16'hEF2C, 16'hD6B2,
 16'hBA6E, 16'hB675, 16'hC6A7, 16'hEC40,
 16'h2ED5, 16'h7818, 16'h7FF9, 16'h7DFA,
 16'h7FFF, 16'h7DEB, 16'h7FFF, 16'h7AEB,
 16'h5110, 16'h11F6, 16'hD602, 16'h9607,
 16'h80EF, 16'h8000, 16'h80D5, 16'h973A,
 16'hC8B8, 16'hFF55, 16'h2B9F, 16'h346B,
 16'h288C, 16'h237D, 16'h237B, 16'h238B,
 16'h2770, 16'h1C94, 16'hF869, 16'hC099,
 16'h8D66, 16'h8199, 16'h8D6A, 16'h9792,
 16'h9D72, 16'hB48A, 16'hD579, 16'hFA85,
 16'h0C7D, 16'hFF82, 16'hDC7D, 16'hC585,
 16'hCD79, 16'hE289, 16'hED74, 16'hDB90,
 16'hC76B, 16'hBC9C, 16'hCD5B, 16'hFCAE,
 16'h3749, 16'h6FC1, 16'h7F35, 16'h7ED3,
 16'h7F26, 16'h67E2, 16'h4516, 16'h1EF1,
 16'h1607, 16'h1D01, 16'h0FF8, 16'hF40F,
 16'hDAEB, 16'hDF1A, 16'hFAE1, 16'h1D23,
 16'h44D9, 16'h622C, 16'h6AD0, 16'h5A34,
 16'h31C7, 16'h153D, 16'h01BF, 16'hF145,
 16'hE6B7, 16'hDB4E, 16'hD6AD, 16'hD158,
 16'hD0A3, 16'hD262, 16'hD498, 16'hDC70,
 16'hE287, 16'hE583, 16'hE973, 16'hD796,
 16'hB662, 16'hAFA6, 16'hC752, 16'hE3B5,
 16'hEC44, 16'hEAC3, 16'hF237, 16'h13CF,
 16'h3E2C, 16'h65D6, 16'h6F2A, 16'h54D5,
 16'h312E, 16'h1FCE, 16'h2A36, 16'h2DC5,
 16'h1E42, 16'h00B5, 16'hE455, 16'hC19F,
 16'hB26F, 16'hB082, 16'hC78E, 16'hF461,
 16'h0FB0, 16'h233F, 16'h3ED3, 16'h681B,
 16'h7EF7, 16'h7EF7, 16'h7F1A, 16'h7ED5,
 16'h543C, 16'h12B3, 16'hD95D, 16'hB894,
 16'hB97A, 16'hC279, 16'hD793, 16'hFC62,
 16'h27A9, 16'h4C4D, 16'h4FBB, 16'h3B3E,
 16'h28C8, 16'h1933, 16'h01D3, 16'hD127,
 16'h9BDE, 16'h8001, 16'h80E8, 16'h8000,
 16'h8DED, 16'hC512, 16'hF8EE, 16'h1E14,
 16'h2BE9, 16'h191A, 16'hF7E2, 16'hD623,
 16'hABD7, 16'h922F, 16'h98CB, 16'hA43C,
 16'h9FBB, 16'h8B4F, 16'h80A6, 16'h8000,
 16'h808B, 16'h9783, 16'hBD6E, 16'hF3A2,
 16'h2D4E, 16'h48C3, 16'h582B, 16'h5DE7,
 16'h5008, 16'h4908, 16'h52EA, 16'h6122,
 16'h74D3, 16'h7F37, 16'h7EC1, 16'h7C46,
 16'h64B5, 16'h404C, 16'h0FB5, 16'hEF48,
 16'hC6BD, 16'h8F3C, 16'h8000, 16'h8027,
 16'h8000, 16'h8006, 16'h850E, 16'h96DE,
 16'hC837, 16'h0EB4, 16'h5761, 16'h7E8A,
 16'h7F8C, 16'h7E5D, 16'h76B9, 16'h6A33,
 16'h6CDF, 16'h7E12, 16'h7FFB, 16'h65F9,
 16'h3611, 16'hFEE8, 16'hD01B, 16'hADE5,
 16'h9C18, 16'h9BEE, 16'hB40A, 16'hE600,
 16'h2EF3, 16'h741D, 16'h7FD0, 16'h7E45,
 16'h7FA4, 16'h6774, 16'h4A74, 16'h2AA4,
 16'h0145, 16'hDBD0, 16'hC31C, 16'hB4F7,
 16'hC0F7, 16'hF31A, 16'h2AD7, 16'h5D36,
 16'h7EC1, 16'h7F44, 16'h7EB9, 16'h5A48,
 16'h12B8, 16'hD547, 16'hB4BC, 16'hAE3E,
 16'hB9CB, 16'hCF29, 16'hDFE4, 16'hE90E,
 16'hE700, 16'hD4F3, 16'hA51A, 16'h8002,
 16'h8034, 16'h8001, 16'h8048, 16'h8001,
 16'h8054, 16'h8002, 16'h805A, 16'h9AA6,
 16'hB357, 16'hCCAD, 16'hE94D, 16'h1CBC,
 16'h4D39, 16'h66D4, 16'h751C, 16'h6FF5,
 16'h64FA, 16'h6718, 16'h7BD6, 16'h7F3C,
 16'h7EB1, 16'h7F62, 16'h7E8D, 16'h7F83,
 16'h7E6E, 16'h7FA0, 16'h5953, 16'h09B9,
 16'hC73E, 16'h97C8, 16'h8134, 16'h8DCF,
 16'hC02F, 16'hF3D1, 16'h0831, 16'h1DCC,
 16'h3639, 16'h3FBF, 16'h264C, 16'hFDA6,
 16'hCC6B, 16'h9881, 16'h8000, 16'h8057,
 16'h95C0, 16'hA527, 16'hAFF2, 16'hCCF4,
 16'hFB27, 16'h26BD, 16'h3560, 16'h3A82,
 16'h459D, 16'h5344, 16'h5AD9, 16'h590C,
 16'h510E, 16'h3ED9, 16'h283F, 16'h0DAA,
 16'hE46B, 16'hA583, 16'h818C, 16'h8000,
 16'h81A0, 16'h8000, 16'h81A4, 16'h8000,
 16'h949C, 16'hE86D, 16'h1487, 16'h1489,
 16'h0363, 16'hF1B4, 16'hFC33, 16'h1DE8,
 16'h3FFC, 16'h4921, 16'h3FC1, 16'h275D,
 16'h1F85, 16'h3699, 16'h5A4B, 16'h7ECE,
 16'h7F1A, 16'h7EFE, 16'h7EED, 16'h7F24,
 16'h7ECD, 16'h5A3E, 16'h42BC, 16'h3249,
 16'h19B4, 16'hF44A, 16'hDABC, 16'hC63A,
 16'hADD4, 16'hAF1D, 16'hC7F2, 16'hE9FE,
 16'hFD14, 16'hFAD8, 16'hF83D, 16'h01AE,
 16'h1066, 16'h2088, 16'h2E88, 16'h226A,
 16'h05A2, 16'hF355, 16'hD2B1, 16'hBE4C,
 16'hC8B5, 16'hDA4C, 16'hE0B0, 16'hD458,
 16'hBF9D, 16'hAE72, 16'hA17C, 16'hAF97,
 16'hD755, 16'hFAC2, 16'h1025, 16'h2CF5,
 16'h4FEF, 16'h672D, 16'h7BB9, 16'h7F60,
 16'h7E88, 16'h6C8F, 16'h4F5A, 16'h32BB,
 16'h1533, 16'h09DD, 16'h0417, 16'h02F2,
 16'h0E07, 16'h35FD, 16'h6E02, 16'h7FFB,
 16'h7E05, 16'h7FF7, 16'h7E0F, 16'h7FE9,
 16'h4E20, 16'hF4D4, 16'hC03B, 16'hA5B5,
 16'h905C, 16'h8091, 16'h8001, 16'h986A,
 16'hBEA9, 16'hD144, 16'hD8CD, 16'hEA24,
 16'hF6EB, 16'hEA07, 16'hC606, 16'h96ED,
 16'h8020, 16'h8000, 16'h8535, 16'hA6C2,
 16'hB745, 16'hC7B6, 16'hE54F, 16'hF2AD,
 16'hED55, 16'hE4AA, 16'hEA56, 16'hE8AB,
 16'hDB53, 16'hCCB0, 16'hC14C, 16'hA4B9,
 16'h8942, 16'h88C3, 16'h9338, 16'h97CD,
 16'h9F2C, 16'hB8DC, 16'hE91C, 16'h20ED,
 16'h500A, 16'h60FE, 16'h5DFA, 16'h5D0F,
 16'h5CE8, 16'h5E21, 16'h4ED6, 16'h2734,
 16'hF3C2, 16'hD748, 16'hC6AE, 16'hBA5B,
 16'hC79D, 16'hEF6B, 16'h188E, 16'h4078,
 16'h6083, 16'h6C80, 16'h647F, 16'h3C81,
 16'h1E81, 16'h107B, 16'h0A88, 16'h0776,
 16'hF28D, 16'hCF6E, 16'hAE98, 16'hAE60,
 16'hC6AA, 16'hDB4B, 16'hE6C1, 16'hF831,
 16'hFFDD, 16'hF116, 16'hF0F6, 16'hFCFF,
 16'h0B0B, 16'h1EEA, 16'h3721, 16'h3FD4,
 16'h3838, 16'h2DBC, 16'h1D4F, 16'h18A7,
 16'h2E60, 16'h4C9C, 16'h6568, 16'h7E94,
 16'h7F70, 16'h7E8B, 16'h7F7A, 16'h7E83,
 16'h7F7F, 16'h7E80, 16'h7F80, 16'h6681,
 16'h3B7F, 16'h2080, 16'h0981, 16'hE27F,
 16'hCD81, 16'hC27F, 16'hBF81, 16'hAD7F,
 16'h8D81, 16'h8001, 16'h8380, 16'h9C81,
 16'hAE7E, 16'hAE82, 16'h9F7E, 16'h8E83,
 16'h807C, 16'h8885, 16'hA978, 16'hCA8B,
 16'hDF72, 16'hF692, 16'h166A, 16'h2A9A,
 16'h4061, 16'h5DA3, 16'h7659, 16'h78AC,
 16'h6850, 16'h61B2, 16'h5D4C, 16'h42B7,
 16'h2146, 16'h06BD, 16'hDF40, 16'hB8C3,
 16'h913B, 16'h8004, 16'h8C3B, 16'h96C4,
 16'hA43E, 16'hAFBF, 16'hD543, 16'h08BB,
 16'h3848, 16'h64B5, 16'h794E, 16'h67AE,
 16'h4556, 16'h22A6, 16'hF45E, 16'hD69E,
 16'hD266, 16'hD897, 16'hE76C, 16'hF691,
 16'h0170, 16'hFF8F, 16'hD973, 16'hA48A,
 16'h8079, 16'h8000, 16'h807F, 16'h8000,
 16'h8086, 16'h8000, 16'h8091, 16'h8B6A,
 16'hBF9A, 16'hF061, 16'h24A5, 16'h4856,
 16'h61B0, 16'h7E48, 16'h7FBF, 16'h7E3B,
 16'h7FCC, 16'h7E2D, 16'h5ED9, 16'h4521,
 16'h32E4, 16'h1818, 16'h13EC, 16'h1C11,
 16'h2DF0, 16'h3B10, 16'h2DEF, 16'h1813,
 16'h02EA, 16'hE61A, 16'hD2E0, 16'hC628,
 16'hAFCE, 16'h963D, 16'h83B7, 16'h8002,
 16'h899D, 16'hB471, 16'hF481, 16'h228C,
 16'h3C68, 16'h52A4, 16'h4F50, 16'h34BD,
 16'h2336, 16'h1CD6, 16'h151F, 16'h12EB,
 16'h270C, 16'h3EFD, 16'h3AFB, 16'h1F0C,
 16'hFCEE, 16'hD516, 16'hB6E8, 16'hA519,
 16'hA4E7, 16'hC818, 16'h00E9, 16'h2716,
 16'h34EA, 16'h3118, 16'h2CE5, 16'h3C1E,
 16'h45DF, 16'h3B23, 16'h31DC, 16'h2325,
 16'h00D9, 16'hDC2A, 16'hC6D2, 16'hC633,
 16'hB8C7, 16'hB03F, 16'hB8BC, 16'hD749,
 16'hFAB2, 16'h0553, 16'h0EA8, 16'h0B5E,
 16'h019D, 16'hFD67, 16'hF095, 16'hE36E,
 16'hEC91, 16'hFB70, 16'hF790, 16'hE36E,
 16'hC295, 16'h9F68, 16'h889C, 16'h805F,
 16'h8002, 16'h8753, 16'hAAB3, 16'hEA48,
 16'h2DBC, 16'h5040, 16'h53C5, 16'h5035,
 16'h57D3, 16'h6824, 16'h66E4, 16'h4D15,
 16'h27F1, 16'h190B, 16'h1CF7, 16'h2B07,
 16'h3FFB, 16'h4F03, 16'h4EFF, 16'h3AFF,
 16'h0F02, 16'hCEFF, 16'h9300, 16'h8003,
 16'h8000, 16'h8002, 16'h8004, 16'h86FB,
 16'hBA06, 16'hF7F9, 16'h2107, 16'h2DF8,
 16'h3C0A, 16'h4EF5, 16'h4D0C, 16'h3BF3,
 16'h280D, 16'h0EF3, 16'hFB0D, 16'hFCF4,
 16'h020B, 16'h00F7, 16'hEA07, 16'hD4FA,
 16'hD105, 16'hC7FD, 16'hC100, 16'hB704,
 16'hAFF7, 16'hC60F, 16'hF3EA, 16'h271C,
 16'h42DE, 16'h5429, 16'h59D0, 16'h4D37,
 16'h49C1, 16'h3848, 16'h1CB0, 16'hFD57,
 16'hDEA3, 16'hCB62, 16'hCC9B, 16'hED68,
 16'h1E94, 16'h576F, 16'h7490, 16'h706F,
 16'h6694, 16'h4D67, 16'h229F, 16'hF85A,
 16'hE2AE, 16'hD748, 16'hC6C4, 16'hB72E,
 16'hAAE1, 16'hB510, 16'hDBFF, 16'h12F1,
 16'h4520, 16'h6ACF, 16'h7F43, 16'h7BAB,
 16'h5767, 16'h2787, 16'h098A, 16'hF366,
 16'hE7A8, 16'hD14D, 16'hA4BD, 16'h8003,
 16'h80CF, 16'h8002, 16'h80D7, 16'h8002,
 16'h8CD3, 16'hDB32, 16'h1DC7, 16'h4943,
 16'h53B0, 16'h4860, 16'h3F8F, 16'h3A82,
 16'h3B6C, 16'h3AA8, 16'h3841, 16'h2DD8,
 16'h230F, 16'h1909, 16'h04E1, 16'hF133,
 16'hCCB9, 16'h965A, 16'h8001, 16'h807A,
 16'h8000, 16'h808F, 16'h8002, 16'h809A,
 16'hA065, 16'hC699, 16'hE96A, 16'h1D91,
 16'h5C78, 16'h7F7C, 16'h7E92, 16'h7F5E,
 16'h7BB3, 16'h6C3C, 16'h75D6, 16'h7F17,
 16'h7EFD, 16'h7EEE, 16'h6725, 16'h57CB,
 16'h4944, 16'h31AF, 16'h1A5C, 16'h159A,
 16'h196D, 16'h0E8F, 16'h0573, 16'h088E,
 16'h286F, 16'h4895, 16'h5E64, 16'h59A5,
 16'h4052, 16'h2AB9, 16'hFD3A, 16'hD0D3,
 16'hAE1F, 16'hA6F1, 16'h9EFF, 16'h8F11,
 16'h95DF, 16'hA42F, 16'hAEC4, 16'hAE49,
 16'hBCAB, 16'hCF60, 16'hDA96, 16'hD972,
 16'hE289, 16'hEF7A, 16'hF384, 16'h017D,
 16'h0883, 16'h0B7C, 16'h1986, 16'h2B77,
 16'h3F8E, 16'h466C, 16'h2D9A, 16'h055F,
 16'hD4A9, 16'hA74F, 16'h86B9, 16'h853F,
 16'hA3C9, 16'hD12F, 16'h01DA, 16'h151C,
 16'h15ED, 16'h150C, 16'h08FA, 16'h0201,
 16'h0003, 16'hF0F8, 16'hD50E, 16'hBCED,
 16'hAB17, 16'hA3E5, 16'hB01E, 16'hC5E0,
 16'hE523, 16'h0AD9, 16'h312B, 16'h57D2,
 16'h6B31, 16'h59CD, 16'h3534, 16'h18CC,
 16'h1034, 16'h12CC, 16'h0735, 16'hE6CA,
 16'hCD36, 16'hC7CB, 16'hD733, 16'hE6D1,
 16'hED29, 16'hFADD, 16'h0C1E, 16'h0FE8,
 16'h0B12, 16'h06F3, 16'h0B07, 16'h1901,
 16'h20F7, 16'h1D11, 16'h04E7, 16'hDF20,
 16'hAED9, 16'h872E, 16'h82CC, 16'h9F3A,
 16'hC2C0, 16'hED43, 16'h15BB, 16'h2E48,
 16'h36B6, 16'h354B, 16'h2CB4, 16'h1A4B,
 16'h19B8, 16'h2444, 16'h37C1, 16'h4539,
 16'h3ACD, 16'h1A2D, 16'h04D9, 16'hF721,
 16'hECE6, 16'hE512, 16'hD6F5, 16'hD704,
 16'hE704, 16'h08F5, 16'h2711, 16'h36E8,
 16'h241F, 16'h0ADC, 16'hF328, 16'hE6D3,
 16'hED32, 16'hECCB, 16'hE338, 16'hDAC4,
 16'hDB3F, 16'hE6BD, 16'h0147, 16'h23B6,
 16'h4D4D, 16'h5DB1, 16'h584F, 16'h4CB1,
 16'h4D4F, 16'h48B1, 16'h4650, 16'h4CAF,
 16'h4050, 16'h2CB3, 16'h1049, 16'hFFBB,
 16'h0041, 16'h0AC3, 16'h1638, 16'h1ECF,
 16'h3829, 16'h5CE0, 16'h6816, 16'h66F5,
 16'h60FF, 16'h500E, 16'h45E5, 16'h3828,
 16'h18CA, 16'h0044, 16'hFAAF, 16'hF45E,
 16'hF095, 16'hEA77, 16'hE67D, 16'hE090,
 16'hBC64, 16'h8DA6, 16'h8000, 16'h80B7,
 16'h8000, 16'h80C2, 16'h8000, 16'h80C9,
 16'h8000, 16'h80C8, 16'h8000, 16'h8DC1,
 16'hC244, 16'hE9B6, 16'h0F50, 16'h38A8,
 16'h4C62, 16'h5794, 16'h6176, 16'h6B80,
 16'h6A89, 16'h656F, 16'h679A, 16'h6B5C,
 16'h66AE, 16'h5749, 16'h45BF, 16'h2739,
 16'hF7CF, 16'hC12B, 16'h92D9, 16'h8024,
 16'h8000, 16'h801F, 16'h8000, 16'h931A,
 16'hC0E7, 16'hF81A, 16'h2AE3, 16'h5320,
 16'h61DE, 16'h5A25, 16'h45D9, 16'h1D27,
 16'hFAD8, 16'hF32A, 16'hF6D3, 16'h0931,
 16'h12CB, 16'h0C38, 16'h06C6, 16'hEF3B,
 16'hCAC3, 16'hAE3F, 16'hA0C0, 16'h9B41,
 16'hA0BF, 16'hA43F, 16'hA0C3, 16'hA53B,
 16'hB8C7, 16'hE038, 16'h08C9, 16'h3237,
 16'h4FC9, 16'h5E36, 16'h6FCB, 16'h7235,
 16'h61CB, 16'h5035, 16'h3FCC, 16'h2332,
 16'h01D0, 16'hE72F, 16'hCED0, 16'hCB33,
 16'hD4CA, 16'hE538, 16'hF7C5, 16'hF83F,
 16'h00BD, 16'h0F47, 16'h0FB4, 16'h1050,
 16'h0BAD, 16'hF457, 16'hDAA5, 16'hCD5E,
 16'hCE9F, 16'hDF64, 16'hFF9B, 16'h2465,
 16'h369A, 16'h3868, 16'h3697, 16'h2869,
 16'h0F98, 16'h0264, 16'h08A1, 16'h135B,
 16'h20AA, 16'h3F50, 16'h53B6, 16'h4A43,
 16'h30C4, 16'h0B35, 16'hDFD4, 16'hBD22,
 16'hA3E8, 16'h980D, 16'hAFFD, 16'hDEFB,
 16'h070D, 16'h19EB, 16'h231C, 16'h2CDC,
 16'h432C, 16'h4FCD, 16'h433A, 16'h37C0,
 16'h2744, 16'h0EB9, 16'hED49, 16'hDBB8,
 16'hD545, 16'hBEBF, 16'hAE3C, 16'hADCA,
 16'hC330, 16'hDBD6, 16'hE321, 16'hECEA,
 16'hF40B, 16'hF800, 16'h01F4, 16'hFD18,
 16'hF3DC, 16'hFB31, 16'h04C2, 16'h014A,
 16'hE9AB, 16'hCB5F, 16'hAD98, 16'h9371,
 16'h8286, 16'h8381, 16'h9679, 16'hB78B,
 16'hF074, 16'h278C, 16'h4274, 16'h4389,
 16'h3B7C, 16'h407F, 16'h5288, 16'h576F,
 16'h429A, 16'h235D, 16'h18AE, 16'h1F46,
 16'h30C6, 16'h492E, 16'h56DD, 16'h5719,
 16'h44F1, 16'h1906, 16'hDC02, 16'hA0F6,
 16'h8010, 16'h8001, 16'h8018, 16'h8002,
 16'h961F, 16'hC6DF, 16'hFD23, 16'h22DC,
 16'h2E24, 16'h3ADC, 16'h4A24, 16'h45DD,
 16'h3722, 16'h22E0, 16'h0B1D, 16'hFAE5,
 16'h0019, 16'h04EA, 16'h0214, 16'hECED,
 16'hD512, 16'hD0ED, 16'hC816, 16'hC0E7,
 16'hB71C, 16'hAFE0, 16'hC624, 16'hF3D9,
 16'h272A, 16'h42D2, 16'h5433, 16'h59C7,
 16'h4D40, 16'h49B8, 16'h3850, 16'h1CAA,
 16'hFD5B, 16'hDEA0, 16'hCB64, 16'hCC9A,
 16'hED68, 16'h1E96, 16'h576B, 16'h7495,
 16'h706A, 16'h6699, 16'h4D62, 16'h22A4,
 16'hF856, 16'hE2B2, 16'hD743, 16'hC6C9,
 16'hB72A, 16'hAAE4, 16'hB50E, 16'hDC01,
 16'h12EE, 16'h4524, 16'h6ACB, 16'h7F45,
 16'h7BAB, 16'h5765, 16'h278B, 16'h0986,
 16'hF369, 16'hE7A6, 16'hD14D, 16'hA4BF,
 16'h8000, 16'h80D0, 16'h8000, 16'h80D8,
 16'h8000, 16'h8CD5, 16'hDB2F, 16'h1DC9,
 16'h4943, 16'h53AF, 16'h4861, 16'h3F8D,
 16'h3A85, 16'h3B69, 16'h3AAA, 16'h3841,
 16'h2DD4, 16'h2317, 16'h1900, 16'h04E9,
 16'hF12B, 16'hCCC3, 16'h964F, 16'h8001,
 16'h806B, 16'h8005, 16'h8081, 16'h8006,
 16'h8090, 16'hA06A, 16'hC69A, 16'hE965,
 16'h1D98, 16'h5C6E, 16'h7F8A, 16'h7E80,
 16'h7F75, 16'h7B97, 16'h6C5B, 16'h75B5,
 16'h7F3A, 16'h7ED7, 16'h7F19, 16'h66F6,
 16'h57FC, 16'h4911, 16'h31E1, 16'h1A2D,
 16'h15C6, 16'h1947, 16'h0AAD, 16'h025D,
 16'h0A9C, 16'h2868, 16'h4897, 16'h6269,
 16'h5C97, 16'h4368, 16'h279B, 16'hFB60,
 16'hCCA8, 16'hAB4D, 16'hA0BF, 16'h9733,
 16'h88DD, 16'h8C12, 16'h9F01, 16'hA8EB,
 16'hAB29, 16'hB8C3, 16'hCF51, 16'hDA9B,
 16'hD779, 16'hE274, 16'hF19E, 16'hF750,
 16'h07C1, 16'h0F2F, 16'h0FE0, 16'h1E14,
 16'h2DF4, 16'h4206, 16'h45FE, 16'h2701,
 16'hF7FE, 16'hBE05, 16'h8DF3, 16'h8001,
 16'h80D9, 16'h9037, 16'hC6B7, 16'h005D,
 16'h158C, 16'h158E, 16'h1356, 16'h04C7,
 16'hEF1C, 16'hE301, 16'hCAE2, 16'hAE3A,
 16'h92AB, 16'h826E, 16'h827B, 16'hA49B,
 16'hC551, 16'hEFC0, 16'h2332, 16'h53D8,
 16'h7E22, 16'h7FE1, 16'h791F, 16'h4ADC,
 16'h262C, 16'h1AC9, 16'h1945, 16'h0CAB,
 16'hEE67, 16'hD784, 16'hDB92, 16'hF358,
 16'hFCBF, 16'h012A, 16'h0BED, 16'h1EFD,
 16'h1D18, 16'h12D5, 16'h0C3C, 16'h15B4,
 16'h235A, 16'h309B, 16'h2E6E, 16'h148B,
 16'hEA79, 16'hAF85, 16'h837A, 16'h818B,
 16'hA16E, 16'hD09B, 16'h0759, 16'h36B4,
 16'h493F, 16'h3BCE, 16'h2D26, 16'h15E5,
 16'h010F, 16'hFFFD, 16'h0FF8, 16'h2812,
 16'h3BE5, 16'h4023, 16'h27D7, 16'h152C,
 16'h0AD4, 16'h012A, 16'hEED9, 16'hCB24,
 16'hB6DF, 16'hBF1D, 16'hDFE9, 16'h0710,
 16'h1EF8, 16'h18FE, 16'h000D, 16'hE2E8,
 16'hD523, 16'hDED3, 16'hE935, 16'hE9C3,
 16'hF144, 16'hF2B7, 16'hF74D, 16'h12B0,
 16'h4651, 16'h7BAE, 16'h7F52, 16'h7EB0,
 16'h7F4D, 16'h78B7, 16'h6B44, 16'h5DC1,
 16'h573A, 16'h3FCA, 16'h2433, 16'hFFD1,
 16'hE92B, 16'hEED8, 16'hF425, 16'hF3DD,
 16'hF123, 16'h00DC, 16'h2426, 16'h31D7,
 16'h352D, 16'h30CE, 16'h1938, 16'h04C1,
 16'hF446, 16'hDBB2, 16'hD158, 16'hD89D,
 16'hE76D, 16'hF789, 16'h0280, 16'h0478,
 16'hF78F, 16'hC76B, 16'h8C9A, 16'h8002,
 16'h80A1, 16'h8001, 16'h80A3, 16'h8001,
 16'h809E, 16'h8001, 16'h8092, 16'h8002,
 16'h8082, 16'hB488, 16'hF76D, 16'h269D,
 16'h5458, 16'h6AB5, 16'h683F, 16'h60CD,
 16'h6226, 16'h5DE6, 16'h5A0F, 16'h6AFB,
 16'h7BFC, 16'h7F0D, 16'h7EEB, 16'h7F1B,
 16'h71E0, 16'h3B23, 16'hF3DC, 16'hAE25,
 16'h8001, 16'h8026, 16'h8002, 16'h8020,
 16'h8005, 16'h801A, 16'hA3E8, 16'hDC18,
 16'h1CE8, 16'h5816, 16'h74EB, 16'h7016,
 16'h4FEA, 16'h2817, 16'h14E6, 16'h1F1D,
 16'h36E0, 16'h3725, 16'h23D5, 16'h1331,
 16'h0AC9, 16'h053F, 16'hF0B8, 16'hEA50,
 16'hF6A8, 16'h135F, 16'h279C, 16'h1F69,
 16'h0E92, 16'h0572, 16'h158A, 16'h3179,
 16'h4986, 16'h587A, 16'h5D88, 16'h5074,
 16'h2692, 16'hFB66, 16'hE2A3, 16'hCF53,
 16'hAAB9, 16'h823A, 16'h8003, 16'h801E,
 16'h8003, 16'h8003, 16'h800A, 16'h8000,
 16'h8C24, 16'hCCD0, 16'h213D, 16'h67B7,
 16'h7F52, 16'h7EA6, 16'h7F60, 16'h6F9D,
 16'h7064, 16'h7E9C, 16'h7F62, 16'h7EA2,
 16'h7F59, 16'h6AAD, 16'h314C, 16'hF7BD,
 16'hC738, 16'hAED4, 16'hAF1F, 16'hD0EF,
 16'h0B04, 16'h4607, 16'h75ED, 16'h7F1F,
 16'h79D7, 16'h5D34, 16'h34BF, 16'h014D,
 16'hCAA8, 16'h9762, 16'h8000, 16'h806F,
 16'h8000, 16'h9877, 16'hBC87, 16'hEF7A,
 16'h2786, 16'h547A, 16'h6B87, 16'h6277,
 16'h4C8C, 16'h3C70, 16'h3494, 16'h3168,
 16'h269C, 16'h0960, 16'hD6A5, 16'h9D55,
 16'h8001, 16'h8048, 16'h8002, 16'h803D,
 16'h8001, 16'h9334, 16'hD0D1, 16'h0C29,
 16'h3ADC, 16'h4620, 16'h36E3, 16'h281B,
 16'h20E6, 16'h0F19, 16'hF3E8, 16'hE718,
 16'hD0E7, 16'hC71A, 16'hD0E4, 16'hEA1F,
 16'h08DE, 16'h1525, 16'h04D7, 16'hE02E,
 16'hBECB, 16'h9D3E, 16'h96B9, 16'hAF50,
 16'hCCA6, 16'hE763, 16'hF395, 16'h0574,
 16'h2083, 16'h5486, 16'h7E71, 16'h7F96,
 16'h7E65, 16'h7F9F, 16'h7E5E, 16'h57A5,
 16'h3E57, 16'h35AC, 16'h2253, 16'h28AC,
 16'h3E56, 16'h57A6, 16'h6061, 16'h4F96,
 16'h3475, 16'h277F, 16'h188E, 16'hF464,
 16'hC7AC, 16'hA743, 16'h9AD0, 16'hAE1B,
 16'hCAFB, 16'hE9EF, 16'hFB28, 16'hE9BF,
 16'hC65A, 16'h968D, 16'h808E, 16'h8000,
 16'h80C2, 16'h8000, 16'h80F1, 16'h81FC,
 16'h8A15, 16'h9BDC, 16'hB430, 16'hC5C6,
 16'hDC42, 16'hFFB9, 16'h3649, 16'h77B8,
 16'h7FFE, 16'h7DC2, 16'h7FFF, 16'h6ED8,
 16'h5819, 16'h4BF9, 16'h40F4, 16'h4220,
 16'h50CA, 16'h594D, 16'h4A9A, 16'h2280,
 16'h0266, 16'hEEB4, 16'hD934, 16'hBEE1,
 16'hB30C, 16'hBF05, 16'hDBED, 16'hE91F,
 16'hE2D6, 16'hC632, 16'hA8CA, 16'h9638,
 16'h81C8, 16'h8534, 16'hA4D2, 16'hC827,
 16'hE9E3, 16'h1011, 16'h1EFC, 16'h18F6,
 16'h0919, 16'hFCD7, 16'h053B, 16'h20B3,
 16'h4D5E, 16'h6B92, 16'h7A7C, 16'h6677,
 16'h4095, 16'h1E61, 16'hEAA8, 16'hB650,
 16'h87B5, 16'h8002, 16'h80BB, 16'h8001,
 16'h83BA, 16'h9249, 16'hB5B3, 16'hD452,
 16'hE5A7, 16'hEE61, 16'h0796, 16'h3075,
 16'h5E7E, 16'h7E8F, 16'h7664, 16'h52A8,
 16'h2E4E, 16'h14BC, 16'h0139, 16'hF6D1,
 16'h0225, 16'h19E5, 16'h3212, 16'h31F6,
 16'h1903, 16'hF104, 16'hC2F4, 16'hA113,
 16'h95E7, 16'hB01F, 16'hDFDC, 16'h1D28,
 16'h48D4, 16'h4F30, 16'h3ACC, 16'h2338,
 16'h19C3, 16'h0743, 16'hF0B7, 16'hDB4F,
 16'hD4AC, 16'hE958, 16'h12A3, 16'h3863,
 16'h3E97, 16'h356F, 16'h308B, 16'h2E7A,
 16'h2382, 16'h1082, 16'h0F7A, 16'h1689,
 16'h1C75, 16'h2B8D, 16'h2C72, 16'h2E8D,
 16'h3476, 16'h2B86, 16'h1280, 16'hF779,
 16'hE48E, 16'hEA6A, 16'hF6A0, 16'hF455,
 16'hF0B8, 16'hE73A, 16'hF6D4, 16'h0B1E,
 16'h14F0, 16'h1502, 16'h210C, 16'h3AE7,
 16'h5D25, 16'h7BD0, 16'h7F39, 16'h7EBF,
 16'h5748, 16'h12B4, 16'hDF4E, 16'hC0B2,
 16'h9B4B, 16'h8000, 16'h803E, 16'h82CD,
 16'h8927, 16'h88E6, 16'h9D0B, 16'hC704,
 16'hF6EC, 16'h2B26, 16'h48C7, 16'h5D4C,
 16'h61A0, 16'h5A74, 16'h4578, 16'h2B9B,
 16'h0E54, 16'hF1BB, 16'hC538, 16'h87D3,
 16'h8000, 16'h80E2, 16'h8000, 16'h80E7,
 16'h8000, 16'h80E0, 16'h8000, 16'h80CD,
 16'h9A41, 16'hC3B0, 16'hDE60, 16'hF38E,
 16'h0684, 16'h2B69, 16'h52AB, 16'h6B41,
 16'h6FD2, 16'h6C1C, 16'h64F5, 16'h5DFB,
 16'h7913, 16'h7EE1, 16'h7F29, 16'h7ED0,
 16'h7F34, 16'h7EC9, 16'h7F3A, 16'h66C6,
 16'h2137, 16'h00CD, 16'hF42C, 16'hFADE,
 16'hF118, 16'hECF3, 16'hF401, 16'h000A,
 16'h0BED, 16'h001B, 16'hE4DE, 16'hC728,
 16'hA8D3, 16'h8331, 16'h8002, 16'h8036,
 16'h8000, 16'h8235, 16'hA8CE, 16'hD12C,
 16'hDFDC, 16'hD71C, 16'hCCED, 16'hD909,
 16'hF701, 16'h19F5, 16'h3215, 16'h42E2,
 16'h2B25, 16'h12D6, 16'h052E, 16'hF7CF,
 16'hE032, 16'hCACE, 16'hC731, 16'hCED2,
 16'hC729, 16'hBEDE, 16'hCB18, 16'hDBF3,
 16'hFD02, 16'h100B, 16'h19E7, 16'h2128,
 16'h04C8, 16'hE948, 16'hDEAA, 16'hDB62,
 16'hE892, 16'hF77A, 16'h067C, 16'h078B,
 16'h0B6F, 16'h0C95, 16'hFF6A, 16'hE095,
 16'hC26D, 16'hBF8E, 16'hB87A, 16'hB07C,
 16'hB490, 16'hB562, 16'hB4AF, 16'hCD3E,
 16'hEED6, 16'h0715, 16'h0B01, 16'hFFEA,
 16'hF12B, 16'hF0BF, 16'h0C58, 16'h3792,
 16'h5784, 16'h5766, 16'h4DAD, 16'h3A42,
 16'h3CCE, 16'h4825, 16'h49E6, 16'h450F,
 16'h38F9, 16'h3B02, 16'h5902, 16'h7DFD,
 16'h7FFF, 16'h7E05, 16'h7FF3, 16'h6E1A,
 16'h37D7, 16'h003A, 16'hD2B2, 16'hB663,
 16'hAF88, 16'hA88E, 16'hB75B, 16'hDFBC,
 16'h162C, 16'h52EE, 16'h7EF7, 16'h7F24,
 16'h6EC2, 16'h5456, 16'h2293, 16'hE983,
 16'hC669, 16'hB3AA, 16'hA445, 16'hA5C9,
 16'hB92B, 16'hD5DF, 16'hE91A, 16'hDFEA,
 16'hCE14, 16'hBDEC, 16'h9716, 16'h80E6,
 16'h8000, 16'h80D6, 16'h8000, 16'h80BD,
 16'h8001, 16'h829D, 16'hB675, 16'hD778,
 16'hF09C, 16'h0950, 16'h06C4, 16'hFD27,
 16'hE4EE, 16'hCEFE, 16'hC316, 16'hD0D7,
 16'hEA3A, 16'h01B5, 16'h1F5C, 16'h3095,
 16'h3879, 16'h427A, 16'h3C91, 16'h3666,
 16'h31A2, 16'h1856, 16'hF7B1, 16'hDB4A,
 16'hC1BA, 16'hAF44, 16'hABBC, 16'hAE45,
 16'hCBB9, 16'hFC4A, 16'h3BB2, 16'h7853,
 16'h7FA7, 16'h7E60, 16'h7F97, 16'h6072,
 16'h2B85, 16'h0183, 16'hE376, 16'hD091,
 16'hD967, 16'hE6A1, 16'hE357, 16'hCEB0,
 16'hBF4B, 16'hBEBA, 16'hBD41, 16'hB4C4,
 16'hB737, 16'hD0CE, 16'hFB2E, 16'h27D6,
 16'h4326, 16'h3FDE, 16'h1F1D, 16'h08E8,
 16'hFD14, 16'hE9F1, 16'hD90A, 16'hC5FB,
 16'hC2FE, 16'hE00A, 16'h0EEF, 16'h3219,
 16'h45DD, 16'h5A2F, 16'h71C4, 16'h7F4A,
 16'h7EA8, 16'h6764, 16'h4C91, 16'h3C7B,
 16'h3179, 16'h3292, 16'h3064, 16'h2DA4,
 16'h1955, 16'hF4B2, 16'hD448, 16'hB7BC,
 16'h8E42, 16'h80BD, 16'h8000, 16'h80B2,
 16'h8000, 16'h839E, 16'hCA71, 16'h097F,
 16'h2C92, 16'h325C, 16'h2DB6, 16'h2338,
 16'h1CDB, 16'h3111, 16'h4502, 16'h4CEC,
 16'h4925, 16'h3FCC, 16'h3841, 16'h31B5,
 16'h2D51, 16'h2DAC, 16'h4555, 16'h71AD,
 16'h7F4E, 16'h7EBA, 16'h7F3A, 16'h7ED5,
 16'h7F1A, 16'h7EFA, 16'h4FEF, 16'h0929,
 16'hC7BE, 16'h915B, 16'h8000, 16'h878F,
 16'hAA57, 16'hD2C2, 16'hF726, 16'h13F0,
 16'h13FC, 16'hF916, 16'hC4DC, 16'h8A2F,
 16'h8000, 16'h813C, 16'h8000, 16'h813E,
 16'h85C6, 16'h8632, 16'h8BD9, 16'hA61A,
 16'hCBF5, 16'hDFFB, 16'hE816, 16'hFBD7,
 16'h0F3E, 16'h21AD, 16'h3069, 16'h2B80,
 16'h0A96, 16'hF156, 16'hDFBE, 16'hD22E,
 16'hB9E3, 16'h980E, 16'h8301, 16'h8CF1,
 16'hAF1B, 16'hD6D9, 16'h0232, 16'h1EC6,
 16'h353F, 16'h3BBE, 16'h3B44, 16'h2ABA,
 16'h0148, 16'hDFB6, 16'hCD4B, 16'hCCB6,
 16'hD748, 16'hE4BA, 16'hF344, 16'hFCBE,
 16'h0241, 16'h01BF, 16'hF141, 16'hCABF,
 16'h9F42, 16'h88BE, 16'h9140, 16'hB2C1,
 16'hDB40, 16'hF0BF, 16'hEA43, 16'hE2BA,
 16'hEA49, 16'h04B4, 16'h1F50, 16'h20AC,
 16'h1558, 16'h08A4, 16'h0261, 16'h1999,
 16'h3F6E, 16'h598B, 16'h617B, 16'h527F,
 16'h3886, 16'h2376, 16'h158E, 16'h086E,
 16'h0795, 16'h0A69, 16'h1698, 16'h2268,
 16'h4698, 16'h7B69, 16'h7F95, 16'h7E6D,
 16'h7F8F, 16'h7E76, 16'h7585, 16'h5681,
 16'h3278, 16'h088F, 16'hE369, 16'hC7A0,
 16'hB356, 16'hB8B5, 16'hDB40, 16'h08CA,
 16'h352E, 16'h57D9, 16'h6721, 16'h60E5,
 16'h3B13, 16'hF6F6, 16'hB703, 16'h8D03,
 16'h8001, 16'h800C, 16'h8003, 16'h8014,
 16'h8001, 16'h801C, 16'h8000, 16'h8022,
 16'h8000, 16'h8024, 16'h8000, 16'h9325,
 16'hB4DA, 16'hC127, 16'hC6D8, 16'hD729,
 16'hE6D8, 16'hF727, 16'h0FD9, 16'h2E26,
 16'h49DA, 16'h6128, 16'h61D6, 16'h492C,
 16'h14D1, 16'hE332, 16'hCACC, 16'hB335,
 16'h9CCB, 16'h9635, 16'hA6CB, 16'hB536,
 16'hBCC9, 16'hC137, 16'hCAC9, 16'hE738,
 16'h06C7, 16'h163A, 16'h22C6, 16'h3838,
 16'h49CB, 16'h5731, 16'h66D3, 16'h682B,
 16'h56D7, 16'h3F25, 16'h27DF, 16'h2E1D,
 16'h44E9, 16'h6710, 16'h7EF6, 16'h7F04,
 16'h7F04, 16'h64F4, 16'h2B13, 16'hECE5,
 16'hBD24, 16'hA3D2, 16'hAF39, 16'hD1BC,
 16'h054E, 16'h2AA8, 16'h2B63, 16'h2D92,
 16'h3179, 16'h307B, 16'h1991, 16'hF064,
 16'hD9A6, 16'hD651, 16'hE5B7, 16'hFC42,
 16'h07C5, 16'h0034, 16'hDCD1, 16'hB82B,
 16'hA1D8, 16'h8E27, 16'h8FD8, 16'hAD2A,
 16'hD2D3, 16'hF331, 16'h05CB, 16'h143A,
 16'h23BE, 16'h484C, 16'h72AA, 16'h7E61,
 16'h7F93, 16'h7E79, 16'h7F7A, 16'h7E94,
 16'h7F5D, 16'h7EB2, 16'h583F, 16'h15D0,
 16'hD722, 16'h9EEB, 16'h8008, 16'h8006,
 16'h8000, 16'h8D20, 16'hAED5, 16'hDB35,
 16'h0EC3, 16'h4042, 16'h67BA, 16'h7F4A,
 16'h7EB4, 16'h5A4D, 16'h22B2, 16'hF74C,
 16'hE4B8, 16'hE744, 16'hF3C1, 16'hF13A,
 16'hE2CB, 16'hD92E, 16'hC6DA, 16'hA91D,
 16'h90ED, 16'h820A, 16'h8EFF, 16'hB4F9,
 16'hEA0D, 16'h19EE, 16'h2717, 16'h1CE6,
 16'h091C, 16'h04E3, 16'h101D, 16'h12E4,
 16'h0F1A, 16'h0BE9, 16'h0213, 16'hFAF3,
 16'h0205, 16'h1504, 16'h27F2, 16'h3718,
 16'h3EDF, 16'h3C2A, 16'h20CC, 16'hE93D,
 16'hC0BB, 16'hAB4D, 16'hADAC, 16'hC359,
 16'hDAA4, 16'hF75D, 16'h08A4, 16'h1058,
 16'h12AE, 16'h0F4B, 16'hF0BE, 16'hCF36,
 16'hB6D7, 16'h971B, 16'h8CF6, 16'h96F6,
 16'hAB20, 16'hB4C8, 16'hBF51, 16'hCA97,
 16'hC780, 16'hBC69, 16'hB3AE, 16'hAE3B,
 16'hB7DB, 16'hD810, 16'hFC02, 16'h18EF,
 16'h221D, 16'h26DA, 16'h2F2D, 16'h36CE,
 16'h5934, 16'h7DCC, 16'h7FFE, 16'h7DD4,
 16'h7FFF, 16'h7DE6, 16'h700F, 16'h5FFF,
 16'h3BF0, 16'h1223, 16'hEDC8, 16'hD84E,
 16'hD99D, 16'hDB77, 16'hE975, 16'hF3A0,
 16'hF84B, 16'h01C9, 16'h0225, 16'h01EB,
 16'h0207, 16'hF106, 16'hDBEE, 16'hC71D,
 16'hCADA, 16'hE02D, 16'hFACF, 16'h0F33,
 16'h18CC, 16'h0933, 16'hDFCF, 16'hAF2F,
 16'h8001, 16'h8026, 16'h8003, 16'h801A,
 16'h9AEC, 16'hB710, 16'hD0F3, 16'hE50A,
 16'hE6F9, 16'hD703, 16'hCF01, 16'hDBFC,
 16'hF306, 16'hFAF8, 16'hF408, 16'hDBFA,
 16'hC804, 16'hCAFE, 16'hE2FF, 16'h0904,
 16'h2AF8, 16'h450E, 16'h59EB, 16'h571C,
 16'h36DD, 16'h152A, 16'h01CE, 16'hEF3B,
 16'hD6BD, 16'hC64A, 16'hC2AF, 16'hC758,
 16'hBEA1, 16'hBA66, 16'hBC94, 16'hB371,
 16'hA68B, 16'h9777, 16'h9E8A, 16'hBD73,
 16'hE991, 16'h136A, 16'h1E9B, 16'h1A60,
 16'h12A6, 16'h1653, 16'h26B6, 16'h2B40,
 16'h2ACA, 16'h232B, 16'h26E1, 16'h3F13,
 16'h61FA, 16'h78F8, 16'h7F16, 16'h7EDD,
 16'h6F2F, 16'h52C5, 16'h3146, 16'h14B1,
 16'h0B57, 16'h1CA3, 16'h3260, 16'h369D,
 16'h3866, 16'h4599, 16'h4566, 16'h379C,
 16'h2860, 16'h20A6, 16'h1553, 16'hFCB4,
 16'hDB44, 16'hB4C5, 16'h9B32, 16'h9CD7,
 16'hA720, 16'hA8E9, 16'hB70F, 16'hCEF8,
 16'hF401, 16'h1505, 16'h15F7, 16'h0B0C,
 16'hFAF2, 16'hE30E, 16'hDAF3, 16'hE30B,
 16'hF2F8, 16'h0904, 16'h1A02, 16'h20F7,
 16'h1A11, 16'h0BE5, 16'h0126, 16'h01D0,
 16'h0C3A, 16'h0BBC, 16'h054D, 16'h12AA,
 16'h2B60, 16'h4996, 16'h5D73, 16'h4E84,
 16'h3C85, 16'h2773, 16'h0294, 16'hDA66,
 16'hB39D, 16'h9563, 16'h809C, 16'h8002,
 16'h8399, 16'h9768, 16'hC796, 16'h006E,
 16'h388D, 16'h5C79, 16'h6281, 16'h5785,
 16'h4074, 16'h2694, 16'h1663, 16'h0FA7,
 16'h074F, 16'hECBA, 16'hCB3E, 16'hAACA,
 16'h8F2D, 16'h81DC, 16'h821B, 16'h97EE,
 16'hCB0A, 16'h04FE, 16'h36F9, 16'h5E10,
 16'h67E7, 16'h5422, 16'h42D7, 16'h322F,
 16'h19CA, 16'h003D, 16'hE9BE, 16'hE747,
 16'hE9B4, 16'hF450, 16'hFAAC, 16'hFB58,
 16'hF0A5, 16'hD15D, 16'hA8A1, 16'h8260,
 16'h8003, 16'h8062, 16'h8003, 16'h8F65,
 16'hAD9A, 16'hC667, 16'hDA98, 16'hF768,
 16'h2399, 16'h5765, 16'h6F9F, 16'h7C5C,
 16'h7EA9, 16'h7952, 16'h6FB3, 16'h7249,
 16'h6EBB, 16'h5740, 16'h49C6, 16'h4533,
 16'h3AD5, 16'h1F24, 16'hFFE2, 16'hE518,
 16'hE6ED, 16'hF10E, 16'hF6F8, 16'hFB03,
 16'h0102, 16'h12F9, 16'h210A, 16'h2CF4,
 16'h310D, 16'h2DF3, 16'h240E, 16'h0BF1,
 16'hE90F, 16'hCEF1, 16'hC10D, 16'hB2F7,
 16'hA406, 16'h9AFD, 16'h90FF, 16'h8705,
 16'h8000, 16'h800A, 16'h8000, 16'h910C,
 16'hBEF4, 16'hF80D, 16'h22F3, 16'h2E0C,
 16'h2DF6, 16'h2406, 16'h26FE, 16'h3EFE,
 16'h5807, 16'h59F4, 16'h5A10, 16'h59EC,
 16'h4618, 16'h3AE4, 16'h2D21, 16'h12D9,
 16'hF82E, 16'hE2CC, 16'hDF38, 16'hE8C5,
 16'hF13D, 16'hFFC3, 16'h0B3C, 16'h08C6,
 16'hFD36, 16'hEECF, 16'hED2C, 16'hF7DA,
 16'hFB1F, 16'hF7E8, 16'hEF10, 16'hECF8,
 16'h0201, 16'h2105, 16'h42F5, 16'h5011,
 16'h42EA, 16'h321A, 16'h15E3, 16'hF31D,
 16'hCEE5, 16'hBF19, 16'hC5EB, 16'hD70F,
 16'hE9F7, 16'hFB01, 16'h070A, 16'hFAEB,
 16'hE022, 16'hC5CE, 16'hAE42, 16'h8BAE,
 16'h8063, 16'h8000, 16'h807F, 16'h8001,
 16'h8098, 16'h965D, 16'hBDAC, 16'hE44C,
 16'hF8BB, 16'h1440, 16'h1DC4, 16'h1E38,
 16'h15CA, 16'h1838, 16'h1AC3, 16'h1844,
 16'h24B1, 16'h275C, 16'h2B98, 16'h3475,
 16'h437D, 16'h5390, 16'h5062, 16'h3FAE,
 16'h3142, 16'h15CE, 16'hFD22, 16'hF2ED,
 16'hE304, 16'hD20B, 16'hC6E8, 16'hBF23,
 16'hB9D4, 16'hBD33, 16'hD0C6, 16'hEA41,
 16'hFFB9, 16'h134C, 16'h2AB0, 16'h3753,
 16'h48AC, 16'h6153, 16'h66AE, 16'h5851,
 16'h4EB1, 16'h4F4D, 16'h49B5, 16'h3F48,
 16'h1EBC, 16'hFB40, 16'hD6C4, 16'hB738,
 16'hA6CB, 16'h9B32, 16'h9ED2, 16'hB72B,
 16'hD8D8, 16'hF324, 16'h00E0, 16'h0B1D,
 16'h12E6, 16'h0F17, 16'h0AEC, 16'h0911,
 16'h08F3, 16'h0108, 16'h00FD, 16'h01FF,
 16'h0005, 16'h08F7, 16'h240C, 16'h44F1,
 16'h6212, 16'h7BED, 16'h7F13, 16'h75EC,
 16'h5015, 16'h22E9, 16'h011A, 16'hE4E4,
 16'hC81C, 16'hB4E5, 16'hB71A, 16'hBEE7,
 16'hC618, 16'hCEE8, 16'hDF19, 16'hEEE8,
 16'hFB16, 16'hF0EC, 16'hDF11, 16'hD0F2,
 16'hD50C, 16'hE8F6, 16'hF807, 16'h00FD,
 16'hF3FE, 16'hE506, 16'hE2F8, 16'hDB09,
 16'hD4F6, 16'hD90B, 16'hD6F3, 16'hE310,
 16'hFFEE, 16'h1914, 16'h23E9, 16'h1D1A,
 16'h0AE3, 16'hFB1F, 16'hFFE1, 16'h091F,
 16'h0EE1, 16'h191E, 16'h19E3, 16'h131B,
 16'h12E8, 16'h2116, 16'h30EB, 16'h3B14,
 16'h37ED, 16'h2E11, 16'h2DF2, 16'h280C,
 16'h14F5, 16'hF80B, 16'hE2F4, 16'hD20E,
 16'hCCF0, 16'hC813, 16'hD1E8, 16'hE91D,
 16'hF7DE, 16'h0928, 16'h12D1, 16'h1036,
 16'h04C0, 16'h014D, 16'hECA6, 16'hDB66,
 16'hDA8E, 16'hE07E, 16'hE976, 16'hED97,
 16'hEC5B, 16'hDBB2, 16'hC644, 16'hB5C5,
 16'hAD31, 16'hB0D9, 16'hCE1E, 16'hF3EA,
 16'h1211, 16'h28F1, 16'h2D0E, 16'h2BF1,
 16'h3013, 16'h38E8, 16'h441E, 16'h40D9,
 16'h4231, 16'h3BC5, 16'h2747, 16'h16AD,
 16'h0A5E, 16'hEF95, 16'hD179, 16'hB979,
 16'hAA96, 16'hB55B, 16'hC0B3, 16'hD740,
 16'hE8CC, 16'hF128, 16'hF6E4, 16'hFB11,
 16'h06F9, 16'h14FE, 16'h190B, 16'h0EEC,
 16'hFD1D, 16'hFADA, 16'h092E, 16'h0FCA,
 16'h163E, 16'h14BA, 16'hFB4D, 16'hD1AD,
 16'hAB58, 16'h86A2, 16'h8064, 16'h8000,
 16'h876D, 16'hAF90, 16'hCF72, 16'hEE8C,
 16'h0977, 16'h1986, 16'h157C, 16'h0F83,
 16'h157E, 16'h1582, 16'h107C, 16'h0187,
 16'hF176, 16'hE28D, 16'hE06F, 16'hF695,
 16'h1367, 16'h309E, 16'h3F5C, 16'h45A9,
 16'h3C52, 16'h1EB3, 16'h0249, 16'hEEBB,
 16'hE340, 16'hDAC5, 16'hD736, 16'hD8CE,
 16'hDC2F, 16'hD6D4, 16'hD529, 16'hD4DA,
 16'hC622, 16'hB4E0, 16'hA520, 16'h9EE0,
 16'hB520, 16'hD6E1, 16'hF71D, 16'h08E5,
 16'h0B18, 16'h0AED, 16'h150D, 16'h22F9,
 16'h2701, 16'h2B04, 16'h26F8, 16'h2D0D,
 16'h3FEC, 16'h571C, 16'h66DC, 16'h6F2C,
 16'h6FCC, 16'h623C, 16'h48BC, 16'h274C,
 16'h0EAC, 16'h055C, 16'h0E9C, 16'h196A,
 16'h1991, 16'h1F73, 16'h2D8A, 16'h2D79,
 16'h2684, 16'h1F7E, 16'h1C82, 16'h1A7C,
 16'h0F87, 16'hF877, 16'hD88B, 16'hBD73,
 16'hB48F, 16'hB76E, 16'hB695, 16'hBF69,
 16'hCE99, 16'hEA64, 16'h06A0, 16'h025C,
 16'hF7A8, 16'hEA55, 16'hD6AD, 16'hD552,
 16'hE2AF, 16'hF750, 16'h0BB1, 16'h1F4F,
 16'h23B1, 16'h1A4F, 16'h0FB0, 16'h0551,
 16'h06AE, 16'h0C53, 16'h08AD, 16'h0153,
 16'h0AAC, 16'h2155, 16'h3BAA, 16'h4957,
 16'h3BA8, 16'h2759, 16'h14A6, 16'hF35C,
 16'hD0A3, 16'hB05D, 16'h97A3, 16'h8C5C,
 16'h88A6, 16'h9358, 16'hAAAB, 16'hD752,
 16'h0BB1, 16'h3F4B, 16'h5DBA, 16'h6240,
 16'h59C6, 16'h4535, 16'h30CF, 16'h1F2D,
 16'h18D8, 16'h0C21, 16'hF2E6, 16'hD514,
 16'hB2F2, 16'h9807, 16'h8D01, 16'h8BF6,
 16'hA114, 16'hD0E4, 16'h0722, 16'h36D8,
 16'h5A2E, 16'h64CD, 16'h4F38, 16'h3FC2,
 16'h3144, 16'h18B6, 16'hFD50, 16'hE8AB,
 16'hE559, 16'hE8A3, 16'hF361, 16'hF69D,
 16'hFD64, 16'hF09C, 16'hD163, 16'hAD9E,
 16'h8562, 16'h8002, 16'h8061, 16'h8003,
 16'h8D5F, 16'hADA2, 16'hC65C, 16'hD8A6,
 16'hF758, 16'h23AB, 16'h5752, 16'h6FB0,
 16'h7C4E, 16'h7EB5, 16'h7948, 16'h6FBC,
 16'h723F, 16'h6EC7, 16'h5733, 16'h49D3,
 16'h4527, 16'h3ADE, 16'h1F1E, 16'hFFE6,
 16'hE515, 16'hE6F1, 16'hF108, 16'hF6FE,
 16'hFAFD, 16'h0106, 16'h12F9, 16'h2107,
 16'h2CF8, 16'h310A, 16'h2DF4, 16'h240D,
 16'h0BF4, 16'hE90A, 16'hCEF8, 16'hC107,
 16'hB2FA, 16'hA404, 16'h9AFF, 16'h90FD,
 16'h8707, 16'h8000, 16'h800A, 16'h8003,
 16'h910C, 16'hBEF3, 16'hF80F, 16'h22EF,
 16'h2E12, 16'h2DEF, 16'h240F, 16'h26F4,
 16'h3F07, 16'h57FF, 16'h59FB, 16'h5A0B,
 16'h59EF, 16'h4617, 16'h3AE2, 16'h2D25,
 16'h12D4, 16'hF833, 16'hE2C7, 16'hDF3D,
 16'hE8C0, 16'hF142, 16'hFFBD, 16'h0B43,
 16'h08BE, 16'hFD40, 16'hEEC2, 16'hED3B,
 16'hF7CB, 16'hFB2D, 16'hF7DB, 16'hEF1C,
 16'hECED, 16'h020B, 16'h20FE, 16'h42F7,
 16'h5014, 16'h42E1, 16'h3229, 16'h15CF,
 16'hF338, 16'hCEC2, 16'hBF43, 16'hC5BA,
 16'hD747, 16'hE9BA, 16'hFB42, 16'h08C5,
 16'hFB34, 16'hDFD3, 16'hC623, 16'hAAE8,
 16'h890D, 16'h8000, 16'h8002, 16'h801F,
 16'h8002, 16'h8042, 16'h90AB, 16'hB966,
 16'hE28B, 16'hFD83, 16'h1870, 16'h239C,
 16'h2358, 16'h19B4, 16'h1C41, 16'h1FC7,
 16'h2034, 16'h27D0, 16'h2A2E, 16'h2BD3,
 16'h362C, 16'h45D2, 16'h5633, 16'h4FC8,
 16'h3E3E, 16'h2BBC, 16'h0E4A, 16'hF7AE,
 16'hE85B, 16'hD99D, 16'hC56B, 16'hB38E,
 16'hA379, 16'h9D7E, 16'hA08C, 16'hB96A,
 16'hDE9F, 16'h0058, 16'h1EB1, 16'h3C46,
 16'h4CC4, 16'h5831, 16'h6BD9, 16'h6F1E,
 16'h61EC, 16'h540A, 16'h5301, 16'h4EF2,
 16'h451B, 16'h27D9, 16'h0134, 16'hD4C0,
 16'hAE4B, 16'h95A8, 16'h8366, 16'h8B8E,
 16'hAE7E, 16'hDF76, 16'h0294, 16'h1962,
 16'h27A8, 16'h2A51, 16'h1DB4, 16'h0E47,
 16'h0BBD, 16'h0640, 16'hF8C2, 16'hEE3D,
 16'hE3C3, 16'hD83F, 16'hE3BD, 16'h0848,
 16'h28B2, 16'h4F56, 16'h72A2, 16'h7E66,
 16'h7C92, 16'h6075, 16'h3884, 16'h1E84,
 16'h0774, 16'hE995, 16'hD161, 16'hC6A7,
 16'hC353, 16'hBCB2, 16'hB749, 16'hB9BC,
 16'hC33F, 16'hC5C5, 16'hB939, 16'hADC8,
 16'hAF37, 16'hC6C9, 16'hE737, 16'hFFC9,
 16'h0539, 16'hF2C4, 16'hE53E, 16'hE4BF,
 16'hE345, 16'hE8B8, 16'hF44B, 16'hFAB2,
 16'h0950, 16'h20AF, 16'h2D52, 16'h2CAE,
 16'h1951, 16'h00B0, 16'hF74F, 16'hFAB3,
 16'h004A, 16'h0BBB, 16'h1F3F, 16'h20C7,
 16'h1A33, 16'h1ED3, 16'h2E27, 16'h3FE0,
 16'h4319, 16'h34EE, 16'h270B, 16'h23FB,
 16'h27FF, 16'h2D07, 16'h19F5, 16'h020F,
 16'hE8ED, 16'hD215, 16'hC0EA, 16'hBD17,
 16'hD0EA, 16'hE714, 16'h00ED, 16'h1512,
 16'h22EF, 16'h2810, 16'h31F2, 16'h280B,
 16'h14F9, 16'h0903, 16'h0900, 16'h14FE,
 16'h1003, 16'h01FD, 16'hE703, 16'hCCFD,
 16'hB703, 16'hAAFC, 16'hAE05, 16'hC5FB,
 16'hE905, 16'h0FFB, 16'h2D04, 16'h2DFD,
 16'h2802, 16'h26FF, 16'h1D01, 16'h06FF,
 16'hF301, 16'hE9FE, 16'hE003, 16'hCEFC,
 16'hC105, 16'hB2FA, 16'hA508, 16'h8EF5,
 16'h800F, 16'h8001, 16'h8C1B, 16'hA3DE,
 16'hBF28, 16'hD8D4, 16'hE530, 16'hE8CC,
 16'hF737, 16'h0BC6, 16'h273D, 16'h42C1,
 16'h4640, 16'h3AC0, 16'h3240, 16'h31C1,
 16'h2D3C, 16'h22C8, 16'h0B33, 16'hE6D4,
 16'hC124, 16'hA0E4, 16'h8D14, 16'h8BF4,
 16'h8F03, 16'hA507, 16'hCCEE, 16'hEF1E,
 16'h15D6, 16'h3B35, 16'h5CC1, 16'h6B47,
 16'h6AB2, 16'h6256, 16'h4CA3, 16'h2D64,
 16'h1593, 16'h0F74, 16'h0488, 16'h057B,
 16'h1284, 16'h247B, 16'h3686, 16'h2E77,
 16'h228E, 16'h0F6D, 16'hF699, 16'hDB60,
 16'hC7A6, 16'hCD54, 16'hDFB5, 16'hF741,
 16'h01C8, 16'h012E, 16'hFFDD, 16'h0219,
 16'hFCF1, 16'hEA03, 16'hD109, 16'hB6ED,
 16'h9F1C, 16'h9EDB, 16'hAF2E, 16'hC2C8,
 16'hD544, 16'hE4B0, 16'hFD59, 16'h0EA0,
 16'h1567, 16'h1892, 16'h2476, 16'h2D81,
 16'h3287, 16'h3B73, 16'h3891, 16'h376D,
 16'h4395, 16'h4469, 16'h3C98, 16'h2668,
 16'h0B97, 16'h006D, 16'hEF8D, 16'hE27A,
 16'hD17E, 16'hC78A, 16'hD16E, 16'hDE9B,
 16'hE35C, 16'hE9AD, 16'hFB48, 16'h0FC3,
 16'h2B32, 16'h44DB, 16'h5417, 16'h4CF6,
 16'h2DFE, 16'h070D, 16'hE9EA, 16'hE31E,
 16'hDEDA, 16'hD22E, 16'hD0CB, 16'hCD3B,
 16'hBCC0, 16'hAF44, 16'hA3B9, 16'hA548,
 16'hB9B9, 16'hDF44, 16'h04C1, 16'h2139,
 16'h31CC, 16'h282F, 16'h1ED6, 16'h1525,
 16'h0FE2, 16'h0B16, 16'hFAF1, 16'hE908,
 16'hDFFF, 16'hE2FB, 16'hE50B, 16'hE4EF,
 16'hD517, 16'hBCE5, 16'hA51D, 16'h90E1,
 16'h8C20, 16'h90E0, 16'h9821, 16'hADDF,
 16'hC81F, 16'hDEE2, 16'hF71D, 16'h15E5,
 16'h3818, 16'h53EC, 16'h650F, 16'h66F7,
 16'h6103, 16'h6803, 16'h79F7, 16'h7F0E,
 16'h79EE, 16'h6516, 16'h52E6, 16'h401E,
 16'h2ADE, 16'h1626, 16'h04D5, 16'h0B30,
 16'h15CC, 16'h1338, 16'h0EC4, 16'h133F,
 16'h0FBF, 16'h0543, 16'hF6BC, 16'hF143,
 16'hECBE, 16'hDF41, 16'hC6C0, 16'hA93E,
 16'h96C5, 16'h9337, 16'h9ACE, 16'hA72B,
 16'hBCDD, 16'hCB1B, 16'hDAED, 16'hE90B,
 16'hE9FD, 16'hE6F9, 16'hE714, 16'hF3DF,
 16'h0B2D, 16'h20C7, 16'h2743, 16'h1EB4,
 16'h1A56, 16'h18A1, 16'h1667, 16'h1291,
 16'h0175, 16'hF087, 16'hE07C, 16'hD082,
 16'hC87F, 16'hC082, 16'hB97B, 16'hAE8B,
 16'hA76D, 16'hAA9B, 16'hAF5D, 16'hBEAD,
 16'hDB49, 16'hFFC2, 16'h1031, 16'h19DC,
 16'h2319, 16'h2DF2, 16'h4A03, 16'h6207,
 16'h66F0, 16'h5D18, 16'h4EE2, 16'h4924,
 16'h4ED6, 16'h462E, 16'h31CF, 16'h1934,
 16'h0BCB, 16'h0234, 16'hF2CD, 16'hEA31,
 16'hECD3, 16'hFB27, 16'h0FE0, 16'h2418,
 16'h34F2, 16'h3B04, 16'h2E06, 16'h15EF,
 16'hFD1B, 16'hF0DE, 16'hDF28, 16'hC6D2,
 16'hAE35, 16'h95C3, 16'h8C44, 16'h95B7,
 16'hA14C, 16'hB4B3, 16'hCF4D, 16'hDFB3,
 16'hF44D, 16'h00B4, 16'h014A, 16'h00B9,
 16'h0743, 16'h0AC3, 16'h0C36, 16'h15D1,
 16'h1A27, 16'h1EE2, 16'h2B16, 16'h36F1,
 16'h3108, 16'h22FE, 16'h0EFC, 16'h020B,
 16'hFFEE, 16'hFB18, 16'h04E2, 16'h0F23,
 16'h0FDB, 16'h0727, 16'hF3D8, 16'hE028,
 16'hD0D7, 16'hC62A, 16'hC0D8, 16'hC725,
 16'hDADE, 16'hF41D, 16'h0BE8, 16'h2314,
 16'h2CF2, 16'h2D05, 16'h2403, 16'h14F5,
 16'h1613, 16'h1EE7, 16'h311F, 16'h3FDA,
 16'h3F2C, 16'h2CCF, 16'h0935, 16'hE9C8,
 16'hCF3A, 16'hB9C5, 16'hB53B, 16'hC2C7,
 16'hE035, 16'h01D0, 16'h192A, 16'h22DD,
 16'h1D1D, 16'h18E9, 16'h1610, 16'h06F8,
 16'hE9FE, 16'hD20D, 16'hCCE8, 16'hD222,
 16'hDED5, 16'hE533, 16'hDFC5, 16'hDF43,
 16'hDAB5, 16'hC752, 16'hB4A9, 16'hA75B,
 16'hA8A3, 16'hBF5C, 16'hDAA7, 16'hED56,
 16'hF2AE, 16'hF44D, 16'hFFB8, 16'h1041,
 16'h23C8, 16'h322F, 16'h3FDB, 16'h461A,
 16'h42F0, 16'h3B06, 16'h2D05, 16'h1EF0,
 16'h051B, 16'hE6DB, 16'hD12D, 16'hBCCD,
 16'hA537, 16'h8EC7, 16'h893A, 16'h8BC6,
 16'h9838, 16'hBCCC, 16'hEA2F, 16'h19D6,
 16'h3824, 16'h3FE3, 16'h3815, 16'h31F4,
 16'h3701, 16'h400B, 16'h48EA, 16'h4620,
 16'h30D7, 16'h1A31, 16'h0BC8, 16'h013E,
 16'hFCBD, 16'h0547, 16'h14B6, 16'h234C,
 16'h2DB3, 16'h244B, 16'h1EB9, 16'h1D42,
 16'h1EC5, 16'h2133, 16'h1ED5, 16'h1F20,
 16'h12ED, 16'hFB07, 16'hE904, 16'hDEF0,
 16'hDC1C, 16'hDED8, 16'hDB34, 16'hCEC1,
 16'hCD49, 16'hD6AF, 16'hD257, 16'hD0A3,
 16'hD263, 16'hD099, 16'hD16A, 16'hD694,
 16'hD76C, 16'hD695, 16'hDF6A, 16'hE998,
 16'hF764, 16'h06A1, 16'h1059, 16'h18AE,
 16'h274B, 16'h37BC, 16'h3B3D, 16'h37CA,
 16'h352F, 16'h36D7, 16'h3B24, 16'h3AE1,
 16'h371B, 16'h30E9, 16'h2B12, 16'h14F2,
 16'hF70A, 16'hE2FA, 16'hCB03, 16'hB000,
 16'hA0FC, 16'hA107, 16'hB2F6, 16'hD10E,
 16'hEEEF, 16'h0214, 16'h08E8, 16'h021C,
 16'hFAE0, 16'hEF25, 16'hE2D5, 16'hE931,
 16'hECCA, 16'hED3B, 16'hECC0, 16'hEA45,
 16'hE4B4, 16'hE754, 16'hE8A5, 16'hE361,
 16'hDB9A, 16'hD569, 16'hDA95, 16'hF16D,
 16'h0B91, 16'h1070, 16'h1490, 16'h0C6E,
 16'hFF97, 16'hFB63, 16'hFCA3, 16'h0B56,
 16'h20B2, 16'h2846, 16'h22C4, 16'h1F30,
 16'h20DC, 16'h2417, 16'h22F7, 16'h18FB,
 16'h0913, 16'hFFDF, 16'hF32D, 16'hE9C8,
 16'hDF42, 16'hD4B4, 16'hCD57, 16'hC69D,
 16'hCD6E, 16'hDA89, 16'hF47F, 16'h147A,
 16'h2E8C, 16'h376E, 16'h2B98, 16'h1264,
 16'hF89F, 16'hE45E, 16'hD2A5, 16'hD858,
 16'hDCAC, 16'hE451, 16'hF8B1, 16'h064D,
 16'h09B4, 16'h004C, 16'hF3B5, 16'hEE4B,
 16'hE9B3, 16'hDB4F, 16'hD7AE, 16'hDA56,
 16'hDFA7, 16'hE65C, 16'hEFA1, 16'hF262,
 16'hF89A, 16'hFC6C, 16'hFB8C, 16'hFF7D,
 16'hF87B, 16'hF08D, 16'hE36A, 16'hDA9E,
 16'hD25A, 16'hD8AF, 16'hEF48, 16'h0BC1,
 16'h2436, 16'h30D3, 16'h2E25, 16'h27E2,
 16'h1D18, 16'h0EED, 16'h050F, 16'hF2F4,
 16'hE70B, 16'hD4F4, 16'hCB0E, 16'hC6F0,
 16'hC711, 16'hCAEE, 16'hD914, 16'hF6E9,
 16'h151B, 16'h3AE0, 16'h5825, 16'h66D7,
 16'h612D, 16'h4CCF, 16'h4035, 16'h30C7,
 16'h1D3C, 16'h06C3, 16'hF83D, 16'hF7C4,
 16'hF73A, 16'hF6C8, 16'hEA37, 16'hDFCB,
 16'hD531, 16'hCAD4, 16'hBA26, 16'hAFE1,
 16'hB919, 16'hCCEC, 16'hE90F, 16'hFAF6,
 16'h0105, 16'hFD01, 16'hF6F9, 16'hF30C,
 16'hFCF0, 16'h0913, 16'h15EB, 16'h2416,
 16'h2DEA, 16'h3116, 16'h2CEA, 16'h2E16,
 16'h37E8, 16'h461A, 16'h52E6, 16'h581A,
 16'h56E5, 16'h461A, 16'h2CE7, 16'h1919,
 16'h04E7, 16'hF819, 16'hE4E6, 16'hCB1B,
 16'hBEE4, 16'hBF1D, 16'hBCE2, 16'hC720,
 16'hD8DD, 16'hE925, 16'hEEDA, 16'hEA26,
 16'hE9DB, 16'hF124, 16'h00DD, 16'h0C22,
 16'h12DF, 16'h0B1E, 16'hFCE7, 16'hF114,
 16'hECF3, 16'hEA05, 16'hEF02, 16'hF2F7,
 16'hF311, 16'hF7E7, 16'hF723, 16'hF2D2,
 16'hEA39, 16'hE4BC, 16'hE04E, 16'hECA9,
 16'h0260, 16'h1899, 16'h2E6D, 16'h378D,
 16'h2779, 16'h1581, 16'h0F85, 16'hFF77,
 16'hF48B, 16'hE675, 16'hDB8A, 16'hDE78,
 16'hEA85, 16'h007F, 16'h157A, 16'h198F,
 16'h1368, 16'h0EA1, 16'h0056, 16'hECB3,
 16'hD743, 16'hC6C6, 16'hC132, 16'hC5D7,
 16'hD120, 16'hDBE9, 16'hED0C, 16'h04FF,
 16'h0EF8, 16'h0F11, 16'h04E6, 16'h0022,
 16'hFFD7, 16'hF32F, 16'hF3CD, 16'hEF36,
 16'hE9C7, 16'hE33B, 16'hD6C4, 16'hD13D,
 16'hCAC3, 16'hCF3B, 16'hE2C8, 16'hFB34,
 16'h15D1, 16'h2829, 16'h2ADE, 16'h2D1A,
 16'h26EF, 16'h2107, 16'h1D03, 16'h0FF3,
 16'h0118, 16'hF2DC, 16'hED30, 16'hE2C4,
 16'hD247, 16'hD0B0, 16'hD158, 16'hD0A0,
 16'hCD67, 16'hC092, 16'hBF77, 16'hC280,
 16'hC887, 16'hD472, 16'hDB95, 16'hDF67,
 16'hDF9C, 16'hDF61, 16'hE09F, 16'hE863,
 16'hFB9B, 16'h0668, 16'h1394, 16'h2270,
 16'h218C, 16'h2278, 16'h1983, 16'h0F83,
 16'h0F76, 16'h1893, 16'h2463, 16'h36A6,
 16'h4351, 16'h3EB8, 16'h373F, 16'h31CA,
 16'h2B2D, 16'h19DC, 16'h071C, 16'hF3EB,
 16'hEF0E, 16'hE6F9, 16'hE501, 16'hEF06,
 16'hF6F3, 16'hFB13, 16'hF0E7, 16'hEA1F,
 16'hE8DC, 16'hEA2A, 16'hE6CF, 16'hE338,
 16'hDEC2, 16'hDC43, 16'hE6BA, 16'hFB48,
 16'h0FB6, 16'h1A4C, 16'h19B1, 16'h1953,
 16'h18AB, 16'h1656, 16'h14A8, 16'h1959,
 16'h20A7, 16'h1A5A, 16'h15A6, 16'h1559,
 16'h14A8, 16'h0F56, 16'h04AE, 16'h004D,
 16'hFFB8, 16'hF744, 16'hE9C0, 16'hDF3C,
 16'hDEC7, 16'hE535, 16'hF2D0, 16'h022C,
 16'h08D8, 16'h0C23, 16'h0FE2, 16'h0B19,
 16'hFCEB, 16'hF112, 16'hE6F0, 16'hE30F,
 16'hDAF3, 16'hD509, 16'hD1FB, 16'hCD02,
 16'hC701, 16'hCAFD, 16'hD703, 16'hDAFD,
 16'hE303, 16'hEEFE, 16'h0101, 16'h0BFF,
 16'h1501, 16'h20FE, 16'h1F03, 16'h19FE,
 16'h1F00, 16'h2302, 16'h1CFB, 16'h1609,
 16'h0FF4, 16'h0910, 16'h04EB, 16'h021B,
 16'h06DE, 16'h102A, 16'h26CD, 16'h3B3D,
 16'h3EB9, 16'h4351, 16'h45A4, 16'h4667,
 16'h448F, 16'h377B, 16'h1C7B, 16'h028E,
 16'hE469, 16'hCFA0, 16'hC658, 16'hCBB0,
 16'hDB49, 16'hEDBC, 16'h0041, 16'h0BC0,
 16'h1240, 16'h0BBF, 16'hFF43, 16'hE3B9,
 16'hD64D, 16'hCFAB, 16'hD05F, 16'hCF96,
 16'hC576, 16'hBD7B, 16'hB997, 16'hC657,
 16'hCEBB, 16'hDC33, 16'hECDF, 16'h020F,
 16'h1303, 16'h19EC, 16'h1F24, 16'h18CC,
 16'h0C45, 16'h06A9, 16'h0168, 16'hFF8A,
 16'hF781, 16'hEC76, 16'hEA91, 16'hE96A,
 16'hF199, 16'hEE66, 16'hE799, 16'hE669,
 16'hDF94, 16'hD870, 16'hD98A, 16'hDA7E,
 16'hD978, 16'hDA93, 16'hE561, 16'hEEAC,
 16'hF446, 16'h0BC7, 16'h162C, 16'h1CE2,
 16'h1D11, 16'h19FC, 16'h14F5, 16'h0918,
 16'h06DD, 16'h052E, 16'h06C8, 16'h0941,
 16'h14B7, 16'h1A4F, 16'h15AD, 16'h0C55,
 16'hFFAB, 16'hF755, 16'hEEAD, 16'hEA4F,
 16'hE8B6, 16'hEF43, 16'hFFC6, 16'h0930,
 16'h0EDC, 16'h1516, 16'h1CF9, 16'h1EF9,
 16'h1915, 16'h15DC, 16'h1632, 16'h15BF,
 16'h0F52, 16'h049E, 16'hF871, 16'hF67F,
 16'hED8F, 16'hEC64, 16'hF8A8, 16'h064E,
 16'h19BA, 16'h233F, 16'h2BC7, 16'h2C35,
 16'h27CD, 16'h1832, 16'h02CE, 16'hEE34,
 16'hD2C8, 16'hC23E, 16'hB7BA, 16'hAF50,
 16'hA7A5, 16'hA666, 16'hB58F, 16'hC27C,
 16'hCD79, 16'hE293, 16'hF460, 16'h06AD,
 16'h1046, 16'h15C6, 16'h102F, 16'h01DC,
 16'h0019, 16'hFCF1, 16'hFD07, 16'hFCFE,
 16'hFD00, 16'hFB01, 16'hEA00, 16'hDEFD,
 16'hDB08, 16'hCCF2, 16'hC115, 16'hB9E2,
 16'hBA28, 16'hBCCD, 16'hC340, 16'hCEB2,
 16'hD95B, 16'hE89A, 16'hF86F, 16'h0489,
 16'h0F7F, 16'h2379, 16'h3190, 16'h3669,
 16'h3B9B, 16'h3663, 16'h319D, 16'h3166,
 16'h3795, 16'h4273, 16'h4581, 16'h3F8D,
 16'h3C64, 16'h3AAC, 16'h3142, 16'h1CD1,
 16'h071B, 16'h00FB, 16'hF3EE, 16'hEA28,
 16'hE2C1, 16'hE556, 16'hEE95, 16'hF87F,
 16'h046E, 16'h0BA3, 16'h0E4E, 16'h07C0,
 16'hFC35, 16'hE3D3, 16'hD827, 16'hD5DE,
 16'hD620, 16'hD2E0, 16'hCC22, 16'hC3D9,
 16'hC02F, 16'hBFC7, 16'hC244, 16'hC7B0,
 16'hD15C, 16'hE598, 16'hFC75, 16'h137D,
 16'h1991, 16'h1960, 16'h12AE, 16'h1047,
 16'h14C3, 16'h1A34, 16'h27D4, 16'h2E25,
 16'h30E1, 16'h271A, 16'h15EA, 16'h0B13,
 16'hF6F1, 16'hE70B, 16'hD6F7, 16'hD108,
 16'hD0F9, 16'hD707, 16'hE2F9, 16'hEA07,
 16'hF2F9, 16'hF406, 16'hF0FC, 16'hF101,
 16'hFB04, 16'hFFF7, 16'h050D, 16'h01F0,
 16'h0112, 16'hFFEC, 16'h0016, 16'h0AE9,
 16'h1918, 16'h22E7, 16'h231A, 16'h26E5,
 16'h241B, 16'h1CE7, 16'h1514, 16'h0FF4,
 16'h0C03, 16'h0906, 16'h00F0, 16'hF719,
 16'hEEDD, 16'hE02F, 16'hD8C5, 16'hD947,
 16'hD0AC, 16'hD25F, 16'hD498, 16'hD771,
 16'hDF87, 16'hEA80, 16'hF27A, 16'hEF8B,
 16'hEC71, 16'hE392, 16'hE46D, 16'hE792,
 16'hEC72, 16'hEF86, 16'hF084, 16'hEF71,
 16'hF39B, 16'hF459, 16'hFAB3, 16'h0540,
 16'h06CE, 16'h1323, 16'h1CED, 16'h2403,
 16'h240B, 16'h26E9, 16'h2721, 16'h23D7,
 16'h212F, 16'h12CC, 16'h0939, 16'h00C3,
 16'hF840, 16'hF6BF, 16'hF73F, 16'hFCC6,
 16'h0134, 16'hFFD3, 16'h0024, 16'hFCE6,
 16'hEF0F, 16'hE6FD, 16'hDFF7, 16'hDF14,
 16'hE8E2, 16'hF128, 16'hF7CE, 16'hFD3C,
 16'hFABB, 16'hF84C, 16'hF3AF, 16'hE955,
 16'hE6A8, 16'hDF5A, 16'hDFA5, 16'hEA5A,
 16'hF6A8, 16'hF855, 16'hFAB0, 16'hF34A,
 16'hE9BD, 16'hED3B, 16'hECCD, 16'hF12B,
 16'hF3DE, 16'hFD19, 16'h01F0, 16'h0106,
 16'h0003, 16'h00F4, 16'h0216, 16'h01E0,
 16'h0028, 16'hFFD1, 16'h0535, 16'h08C6,
 16'h0B3D, 16'h06C2, 16'h023F, 16'h00C1,
 16'h003E, 16'h01C3, 16'h0B3C, 16'h18C7,
 16'h1F34, 16'h20D2, 16'h2127, 16'h19E2,
 16'h0F15, 16'h04F2, 16'hFB07, 16'hF401,
 16'hECF8, 16'hEA0E, 16'hF3EC, 16'h011A,
 16'h04E1, 16'h0924, 16'h0BD6, 16'h102F,
 16'h0BCE, 16'h0234, 16'hFACB, 16'hF435,
 16'hF3CC, 16'hF732, 16'hFCD2, 16'h0028,
 16'hFFDF, 16'hF31A, 16'hE6ED, 16'hDB0C,
 16'hCEFC, 16'hC7FB, 16'hCB0F, 16'hD1E7,
 16'hDC22, 16'hE6D5, 16'hED34, 16'hF7C3,
 16'h0146, 16'h08B2, 16'h0C54, 16'h15A7,
 16'h1D5C, 16'h23A2, 16'h245F, 16'h1CA1,
 16'h135E, 16'h0AA3, 16'h075B, 16'hFCA8,
 16'hF154, 16'hE9B1, 16'hE348, 16'hE4BF,
 16'hE03B, 16'hDECC, 16'hDF2C, 16'hE2DD,
 16'hF118, 16'hF6F3, 16'hFB03, 16'h0107,
 16'h06F0, 16'h0C17, 16'h12E2, 16'h1526,
 16'h0FD2, 16'h0C35, 16'h08C4, 16'h0142,
 16'h01BB, 16'h0746, 16'h0FB8, 16'h1F4B,
 16'h20B2, 16'h1D51, 16'h1CAD, 16'h1353,
 16'h08AE, 16'hFD50, 16'hFAB3, 16'hFB4A,
 16'hF7BA, 16'hFB41, 16'hF7C4, 16'hF438,
 16'hF6CC, 16'hFD30, 16'hFCD5, 16'hFD24,
 16'h00E4, 16'h0014, 16'hFFF4, 16'hFB04,
 16'hF803, 16'hF6F6, 16'hF412, 16'hEEE5,
 16'hF124, 16'hECD3, 16'hEA35, 16'hECC5,
 16'hEF40, 16'hF7BC, 16'h0047, 16'h00B7,
 16'h0149, 16'h04B8, 16'h0747, 16'h0EBA,
 16'h0B45, 16'h0ABC, 16'h0C42, 16'h08C1,
 16'h003B, 16'hFACA, 16'hF731, 16'hF0D4,
 16'hEA27, 16'hE9DD, 16'hE920, 16'hE8E2,
 16'hED1E, 16'hECE2, 16'hF11E, 16'hF6E0,
 16'hFB23, 16'h01D9, 16'h0B2C, 16'h0BCF,
 16'h1036, 16'h0BC5, 16'h0740, 16'h06BB,
 16'h074A, 16'h06B2, 16'h0251, 16'h00AC,
 16'h0056, 16'h01AA, 16'h0056, 16'h00AB,
 16'hFD52, 16'h04B2, 16'h0248, 16'hFCC0,
 16'hFD38, 16'hF6D1, 16'hF326, 16'hF3E3,
 16'hF412, 16'hF6FB, 16'hF6F8, 16'hF315,
 16'hF0DE, 16'hEF2D, 16'hF0CA, 16'hF43E,
 16'hF6BB, 16'hF84B, 16'hF7B0, 16'hF454,
 16'hF3A9, 16'hEF58, 16'hF0A9, 16'hF356,
 16'hF6AC, 16'hF450, 16'hF3B5, 16'hF345,
 16'hF2C2, 16'hF837, 16'hFCCF, 16'h002B,
 16'hFCDB, 16'hFD1F, 16'hFCE7, 16'h0214,
 16'h08EF, 16'h0B0F, 16'h08F2, 16'h070E,
 16'h06F1, 16'h0710, 16'h08EE, 16'h0C15,
 16'h0FE7, 16'h0F1E, 16'h08DB, 16'h022D,
 16'hFCCA, 16'hFB3F, 16'hF6B9, 16'hF34F,
 16'hF2A9, 16'hF45E, 16'hFA9B, 16'hFB6B,
 16'hFF90, 16'hFD75, 16'hF687, 16'hF37C,
 16'hF080, 16'hEF84, 16'hF67A, 16'h0087,
 16'h0879, 16'h0985, 16'h087F, 16'h077D,
 16'h0187, 16'hFB74, 16'hF692, 16'hF867,
 16'hFFA1, 16'h0556, 16'h01B2, 16'h0247,
 16'hFFC0, 16'hF738, 16'hF2D0, 16'hF427,
 16'hF3E2, 16'hF817, 16'hFFF0, 16'h0108,
 16'h04FF, 16'h01FC, 16'h0009, 16'hFCF3,
 16'hF710, 16'hECEE, 16'hE713, 16'hE4EE,
 16'hDF10, 16'hDAF2, 16'hD90C, 16'hDFF7,
 16'hE304, 16'hE903, 16'hF3F5, 16'h0114,
 16'h0AE2, 16'h1028, 16'h14CD, 16'h103F,
 16'h08B5, 16'h0257, 16'hFF9C, 16'hF872,
 16'hF380, 16'hF48F, 16'hEE61, 16'hE9AE,
 16'hE243, 16'hDCCC, 16'hDA27, 16'hD5E5,
 16'hD80F, 16'hDCFC, 16'hE1FA, 16'hEA0E,
 16'hF1ED, 16'hF518, 16'hFEE3, 16'h0620,
 16'h0ADE, 16'h1123, 16'h1BE0, 16'h251A,
 16'h26ED, 16'h280B, 16'h1FFE, 16'h1AF8,
 16'h1814, 16'h19DE, 16'h1E32, 16'h21BD,
 16'h2254, 16'h249B, 16'h2776, 16'h2379,
 16'h1998, 16'h0B56, 16'h08BD, 16'hFD30,
 16'hF2E3, 16'hED0C, 16'hE902, 16'hECF1,
 16'hF31C, 16'hFAD8, 16'hFD33, 16'h01C4,
 16'h0542, 16'hFFBA, 16'hF349, 16'hECB4,
 16'hE94E, 16'hE8B2, 16'hE74C, 16'hE2B8,
 16'hDF42, 16'hDAC5, 16'hD734, 16'hD8D3,
 16'hDB26, 16'hDFE1, 16'hE918, 16'hF6EF,
 16'h000A, 16'h01FD, 16'hFFFC, 16'hFD0B,
 16'hFFF0, 16'h0213, 16'h0BEB, 16'h1917,
 16'h1CE8, 16'h1A19, 16'h15E5, 16'h0F1D,
 16'h0AE1, 16'hFD22, 16'hF0DB, 16'hE727,
 16'hDFD6, 16'hE32D, 16'hE8D0, 16'hEF33,
 16'hF7CA, 16'h003A, 16'h00C0, 16'h0047,
 16'hFFB1, 16'h0258, 16'h01A0, 16'h0567,
 16'h0092, 16'hFD76, 16'hFC83, 16'hFB84,
 16'h0475, 16'h1090, 16'h186E, 16'h1A94,
 16'h1E6A, 16'h1A96, 16'h156C, 16'h0F90,
 16'h0A77, 16'h027F, 16'h018C, 16'hFB68,
 16'hF2A6, 16'hF14A, 16'hE4C7, 16'hDC27,
 16'hDAEC, 16'hD901, 16'hDC11, 16'hDEDE,
 16'hE332, 16'hE9BE, 16'hF353, 16'hF39C,
 16'hF373, 16'hF27F, 16'hEA8D, 16'hEC6B,
 16'hED9A, 16'hF063, 16'hF19E, 16'hF263,
 16'hEF9A, 16'hF26B, 16'hF48E, 16'hF77B,
 16'hFD7B, 16'h0490, 16'h0F64, 16'h15A8,
 16'h1A4C, 16'h1CC0, 16'h2134, 16'h20D9,
 16'h211A, 16'h1EF2, 16'h1304, 16'h0904,
 16'h01F7, 16'hFB0B, 16'hFAF4, 16'hFB0D,
 16'hFFF3, 16'h020D, 16'h00F3, 16'h010B,
 16'hFAFA, 16'hF3FF, 16'hEA09, 16'hE4EE,
 16'hE31C, 16'hE8DB, 16'hF32E, 16'hF6C8,
 16'hFB41, 16'hF7B8, 16'hF84E, 16'hF7AE,
 16'hED54, 16'hE8AA, 16'hE558, 16'hE6A7,
 16'hED58, 16'hF7AB, 16'hFB50, 16'hFCB6,
 16'hF444, 16'hECC3, 16'hED34, 16'hEED5,
 16'hF322, 16'hF6E8, 16'h000E, 16'h01FC,
 16'h00F9, 16'h0012, 16'h00E4, 16'h0226,
 16'h01D1, 16'h0037, 16'h01C2, 16'h0544,
 16'h08B8, 16'h0B4A, 16'h06B4, 16'h024F,
 16'h00AF, 16'h0051, 16'h01B0, 16'h0B4C,
 16'h18BA, 16'h1F3F, 16'h20C8, 16'h2131,
 16'h19D5, 16'h0F25, 16'h04E2, 16'hFB16,
 16'hF3F2, 16'hED05, 16'hEA05, 16'hF3F1,
 16'h0119, 16'h04DE, 16'h0929, 16'h0BD2,
 16'h1031, 16'h0BCD, 16'h0234, 16'hFACB,
 16'hF435, 16'hF3CC, 16'hF733, 16'hFCD0,
 16'h002A, 16'hFFDC, 16'hF31E, 16'hE6EA,
 16'hDB0E, 16'hCEFA, 16'hC7FD, 16'hCB0D,
 16'hD1E9, 16'hDC21, 16'hE6D4, 16'hED37,
 16'hF7C0, 16'h0147, 16'h08B4, 16'h0C50,
 16'h15AB, 16'h1D5A, 16'h23A3, 16'h245F,
 16'h1CA1, 16'h135D, 16'h0AA5, 16'h0759,
 16'hFCAB, 16'hF150, 16'hE9B5, 16'hE346,
 16'hE4C0, 16'hE039, 16'hDECF, 16'hDF28,
 16'hE2E2, 16'hF115, 16'hF6F3, 16'hFB06,
 16'h0100, 16'h06FB, 16'h0C0B, 16'h12EF,
 16'h1517, 16'h0FE1, 16'h0C27, 16'h08D2,
 16'h0135, 16'h01C5, 16'h073F, 16'h0FBD,
 16'h1F47, 16'h20B5, 16'h1D4F, 16'h1CAD,
 16'h1358, 16'h08A3, 16'hFD60, 16'hFA9E,
 16'hFB63, 16'hF79D, 16'hFB63, 16'hF79C,
 16'hF465, 16'hF69B, 16'hFD63, 16'hFCA0,
 16'hFD5C, 16'h00A9, 16'h0051, 16'hFFB6,
 16'hF843, 16'hF6C4, 16'hF434, 16'hF2D5,
 16'hF122, 16'hF2E8, 16'hED0E, 16'hE9FB,
 16'hECFC, 16'hF10E, 16'hF7E9, 16'h0020,
 16'h01D7, 16'h0131, 16'h04C8, 16'h073E,
 16'h0EBF, 16'h0B42, 16'h0ABD, 16'h0944,
 16'h04BB, 16'hFD47, 16'hF7B9, 16'hF345,
 16'hECBE, 16'hE73E, 16'hE6C6, 16'hE737,
 16'hE4CD, 16'hE92E, 16'hE8D7, 16'hEA25,
 16'hF0DE, 16'hF31F, 16'hFAE3, 16'h071D,
 16'h04E3, 16'h091E, 16'h06E0, 16'h0021,
 16'h01DF, 16'h0521, 16'h08DF, 16'h0B21,
 16'h08DF, 16'h0721, 16'h06E0, 16'h021E,
 16'h00E3, 16'hFD1C, 16'h00E7, 16'h0117,
 16'hFFEB, 16'h0011, 16'hFCF3, 16'hFD0B,
 16'hFCF8, 16'hFD03, 16'h0002, 16'h00F8,
 16'h0110, 16'hFCE8, 16'hF41F, 16'hF2D9,
 16'hF42E, 16'hF2CD, 16'hF137, 16'hEEC5,
 16'hE73E, 16'hE8BE, 16'hE747, 16'hE8B3,
 16'hEF53, 16'hF0A8, 16'hF35D, 16'hF39F,
 16'hF464, 16'hF398, 16'hF86D, 16'h048F,
 16'h0576, 16'h0486, 16'h077C, 16'h0681,
 16'h0F84, 16'h1877, 16'h198F, 16'h146A,
 16'h109D, 16'h0F5D, 16'h0BA9, 16'h0852,
 16'h07B2, 16'h0A4B, 16'h09B7, 16'h0048,
 16'hF8B8, 16'hF749, 16'hF4B6, 16'hEE4B,
 16'hE9B3, 16'hE851, 16'hE5A9, 16'hE95F,
 16'hEF97, 16'hF674, 16'hF881, 16'hF68B,
 16'hF369, 16'hF2A2, 16'hF151, 16'hF6BD,
 16'h0035, 16'h04DB, 16'h0515, 16'h00F8,
 16'hFCFC, 16'hF110, 16'hE8E4, 16'hE329,
 16'hE6CA, 16'hF142, 16'hFAB3, 16'h0557,
 16'h04A0, 16'h0268, 16'hFF91, 16'hF475,
 16'hEE88, 16'hEA7A, 16'hE483, 16'hE37E,
 16'hE483, 16'hE97D, 16'hEC84, 16'hEF79,
 16'hF689, 16'hFB76, 16'hFC8D, 16'hFD6F,
 16'h0195, 16'h0166, 16'hFFA0, 16'h005A,
 16'hFFAC, 16'hFD4E, 16'hFCB9, 16'h0140,
 16'h04C7, 16'h0C32, 16'h0FD5, 16'h1524,
 16'h12E3, 16'h0B16, 16'h04F1, 16'hFB08,
 16'hF7FF, 16'hEEF9, 16'hED0F, 16'hE6E9,
 16'hE31E, 16'hE2DC, 16'hE02A, 16'hE2D0,
 16'hE736, 16'hEEC5, 16'hFD3F, 16'h08BD,
 16'h0947, 16'h12B6, 16'h104D, 16'h0FB0,
 16'h0F52, 16'h0FAD, 16'h1354, 16'h12AB,
 16'h1554, 16'h15AF, 16'h0F4F, 16'h06B3,
 16'h0149, 16'hF6BA, 16'hF844, 16'hF3C0,
 16'hF73B, 16'hFFCA, 16'h0730, 16'h0FD7,
 16'h1023, 16'h12E3, 16'h0C16, 16'h0BF1,
 16'h0709, 16'hFCFD, 16'hF7FD, 16'hED09,
 16'hE4F2, 16'hE513, 16'hE9E8, 16'hED1C,
 16'hF2E0, 16'h0026, 16'h04D5, 16'h072E,
 16'h08CF, 16'h0732, 16'h04CE, 16'h0532,
 16'h04CF, 16'h022F, 16'h00D3, 16'hFD2A,
 16'hFFD8, 16'hFB26, 16'hF2DF, 16'hED1B,
 16'hE6EA, 16'hDB10, 16'hD4F6, 16'hCF05,
 16'hD200, 16'hDEFB, 16'hE708, 16'hF0F5,
 16'hF40E, 16'hF3EF, 16'hF415, 16'hF6E7,
 16'hFB1B, 16'h04E5, 16'h011B, 16'h01E4,
 16'h051D, 16'h01E2, 16'h0520, 16'h08DE,
 16'h0B23, 16'h0EDB, 16'h1627, 16'h18D8,
 16'h1D29, 16'h19D5, 16'h132E, 16'h0ACD,
 16'h0538, 16'hFAC4, 16'hF840, 16'hF7BC,
 16'hEF48, 16'hF2B2, 16'hFB55, 16'h00A5,
 16'h0062, 16'h0196, 16'h0172, 16'hFF87,
 16'hF480, 16'hEE79, 16'hE98D, 16'hE86E,
 16'hE797, 16'hE465, 16'hE99E, 16'hE65E,
 16'hE5A5, 16'hE85A, 16'hEFA7, 16'hF658,
 16'hFDA8, 16'h0658, 16'h09A8, 16'h085A,
 16'h02A3, 16'h0160, 16'h009D, 16'hFF65,
 16'h009A, 16'hFF68, 16'hFD95, 16'hFC6E,
 16'hF48E, 16'hF276, 16'hEA88, 16'hE87A,
 16'hEA83, 16'hE87F, 16'hED7F, 16'hEC84,
 16'hF179, 16'hF08A, 16'hF372, 16'hF393,
 16'hFB69, 16'h049A, 16'h0563, 16'h08A0,
 16'h055D, 16'h06A7, 16'h0254, 16'h06B1,
 16'h024A, 16'h04BB, 16'h0B40, 16'h08C5,
 16'h0C35, 16'h08D1, 16'h0929, 16'hFFDD,
 16'hFB1D, 16'hFAE9, 16'hF311, 16'hECF4,
 16'hE908, 16'hECFB, 16'hF102, 16'hFB01,
 16'hFFFC, 16'hFD07, 16'h01F7, 16'h0109,
 16'hFFF8, 16'h0007, 16'hFFFA, 16'h0004,
 16'hFFFE, 16'h0000, 16'hFD03, 16'hFCFB,
 16'hFD05, 16'hFCFB, 16'hFD05, 16'h00FB,
 16'h0206, 16'hFFF7, 16'h000D, 16'hFCEF,
 16'hFD15, 16'h00E8, 16'h0118, 16'h01E9,
 16'h0216, 16'hFFED, 16'h000F, 16'hFCF5,
 16'hF707, 16'hF2FD, 16'hEF00, 16'hEA04,
 16'hECF6, 16'hF411, 16'hF7E8, 16'hFB1E,
 16'h00DD, 16'h0128, 16'hFFD3, 16'hFD31,
 16'hF7CA, 16'hFB3B, 16'hFCC1, 16'h0043,
 16'hFFB8, 16'h004D, 16'hFFAF, 16'hFD53,
 16'h00AE, 16'h024F, 16'h08B5, 16'h0947,
 16'h0ABD, 16'h0C3E, 16'h0AC9, 16'h0B2E,
 16'h06DC, 16'h021A, 16'h01F1, 16'h0002,
 16'hF80B, 16'hF2E8, 16'hF326, 16'hEECD,
 16'hF140, 16'hF3B3, 16'hF459, 16'hFF9C,
 16'h026F, 16'h0088, 16'h0280, 16'h0478,
 16'h0290, 16'h0168, 16'h009F, 16'hFF5C,
 16'hFDA6, 16'hFC5A, 16'hFDA5, 16'hFC5D,
 16'hFDA0, 16'hFA65, 16'hF493, 16'hF377,
 16'hF37D, 16'hF091, 16'hEF61, 16'hF2AC,
 16'hF446, 16'hF7CA, 16'hFB25, 16'hFCEC,
 16'h0003, 16'h010E, 16'h01E2, 16'h052D,
 16'h04C4, 16'h054B, 16'h06A8, 16'h0563,
 16'h0493, 16'h0576, 16'h0683, 16'h0582,
 16'h047A, 16'h078A, 16'h0A74, 16'h098C,
 16'h0675, 16'h0188, 16'hFC7D, 16'hFB7E,
 16'hFC88, 16'hFB71, 16'hFF96, 16'hFD61,
 16'hFFA9, 16'h004E, 16'h00BB, 16'h023B,
 16'h01CE, 16'h0229, 16'hFCE0, 16'hFD18,
 16'hF3EF, 16'hF30A, 16'hF2FD, 16'hF2FD,
 16'hF407, 16'hF0F7, 16'hF30A, 16'hF2F6,
 16'hF30A, 16'hF7F6, 16'h0209, 16'h00F9,
 16'h0205, 16'h00FD, 16'hFD00, 16'h0003,
 16'hF7FA, 16'hF80A, 16'hFFF1, 16'h0013,
 16'hFFE9, 16'hFD1B, 16'h00E2, 16'h0120,
 16'h00E0, 16'hFD1E, 16'hF3E4, 16'hF11A,
 16'hE8E9, 16'hE914, 16'hE8F0, 16'hE70A,
 16'hE9FD, 16'hEEFD, 16'hF409, 16'hFAF1,
 16'h0514, 16'h0AE7, 16'h101F, 16'h0EDC,
 16'h0B29, 16'h04D1, 16'h0034, 16'hFCC8,
 16'hFD3C, 16'hFFC2, 16'h003F, 16'hFFC0,
 16'h0040, 16'hFFC0, 16'hFD40, 16'hFCC2,
 16'hF43A, 16'hF2CA, 16'hF332, 16'hF0D2,
 16'hF12A, 16'hF2DB, 16'hF41E, 16'hF7EA,
 16'hFB0E, 16'hFCF9, 16'h0101, 16'h0105,
 16'hFFF5, 16'h0010, 16'h00EB, 16'h011A,
 16'hFCE2, 16'hFD21, 16'hFCDD, 16'hF425,
 16'hF6D9, 16'hFB28, 16'h00D7, 16'h002A,
 16'hFFD7, 16'h0027, 16'hFFDA, 16'h0026,
 16'hFFDA, 16'h0026, 16'hF7D9, 16'hF829,
 16'hF6D6, 16'hFB2B, 16'h00D3, 16'h002F,
 16'h00CF, 16'h0234, 16'h04C9, 16'h0B39,
 16'h0AC5, 16'h0B3D, 16'h08C0, 16'h0245,
 16'h04B6, 16'h014D, 16'h01B0, 16'hFD52,
 16'hFAAD, 16'hFD55, 16'hFCAA, 16'hF456,
 16'hF2AA, 16'hF855, 16'hFAAD, 16'h0152,
 16'hFFB0, 16'hF84C, 16'hF6B8, 16'hF744,
 16'hF7C1, 16'hFB3A, 16'hF7CB, 16'hFB2F,
 16'hFAD7, 16'hF723, 16'hFAE4, 16'hF714,
 16'hFAF4, 16'h0104, 16'h0005, 16'hFFF2,
 16'h0016, 16'hFFE2, 16'h0026, 16'hFFD3,
 16'hFD33, 16'hFCC8, 16'hFD3D, 16'hFCBE,
 16'hFD46, 16'hFCB7, 16'hFD4B, 16'hF6B5,
 16'hF74A, 16'hFAB7, 16'hFB46, 16'h00C0,
 16'h003A, 16'hFFCC, 16'h002C, 16'hFFDD,
 16'h0019, 16'hFFF3, 16'h0000, 16'h000D,
 16'hFCE6, 16'hFD27, 16'hFCCB, 16'hFD43,
 16'hFCAF, 16'hF85F, 16'hF793, 16'hF87A,
 16'hF67A, 16'hF791, 16'hF765, 16'hFBA4,
 16'h0054, 16'hF8B1, 16'h004D, 16'h00B4,
 16'hF74C, 16'hF8B2, 16'hF651, 16'hF7AB,
 16'hFA5B, 16'hF79C, 16'hFA6F, 16'hF786,
 16'hF785, 16'hFB6F, 16'hF69D, 16'hF857,
 16'hF7B6, 16'hF43D, 16'hF6CF, 16'hF825,
 16'hFAE6, 16'hF810, 16'hFAFA, 16'h00FD,
 16'hF80B, 16'hFAED, 16'hFB1B, 16'hFADE,
 16'h0127, 16'hFFD5, 16'h002E, 16'hFFD0,
 16'h0031, 16'hFFCE, 16'hFD32, 16'hFCCE,
 16'hFD32, 16'hFCCF, 16'hFD30, 16'hFCD0,
 16'hFD31, 16'hFCCE, 16'hFD34, 16'hFCC9,
 16'hF83A, 16'hF7C4, 16'hF73F, 16'hFABD,
 16'h0148, 16'hFFB1, 16'h0057, 16'hFFA2,
 16'h0064, 16'hFF97, 16'hF86E, 16'hF68C,
 16'hFB7B, 16'h007E, 16'h0089, 16'hFF70,
 16'h0095, 16'hFF67, 16'h009C, 16'hFF63,
 16'hF89D, 16'hFF64, 16'h009A, 16'hFF68,
 16'h0095, 16'h0071, 16'h0189, 16'h007E,
 16'h0079, 16'hFC91, 16'hFD66, 16'hFCA5,
 16'hFD4F, 16'hFCBC, 16'h0138, 16'h00D5,
 16'hFD1E, 16'h00F0, 16'hFD01, 16'hFD0D,
 16'hFCE5, 16'hFD29, 16'hFCCA, 16'hFD43,
 16'hFCAF, 16'h0060, 16'hFF92, 16'hF47B,
 16'hF379, 16'hF490, 16'hF36A, 16'hF79C,
 16'h015D, 16'h01A9, 16'hFF52, 16'h00B2,
 16'hFF4C, 16'h00B5, 16'hFF4A, 16'hF4B6,
 16'hF34B, 16'hF8B3, 16'h0052, 16'h00A8,
 16'hFF5E, 16'h009B, 16'hFF6B, 16'h0090,
 16'hF377, 16'hF481, 16'hF388, 16'hF46E,
 16'h019C, 16'h005A, 16'hFFB0, 16'h0047,
 16'hFFC2, 16'h0034, 16'hFFD5, 16'h0022,
 16'hFFE7, 16'hFD00, 16'h11F6, 16'h0103,
 16'h0103, 16'hFFF7, 16'hFD10, 16'hFCEA,
 16'hFD1B, 16'hFCE1, 16'hFD21, 16'h00DE,
 16'h0123, 16'h06DC, 16'h0524, 16'h00DE,
 16'h001E, 16'hFCE7, 16'hF713, 16'hF3F3,
 16'hF708, 16'hFAFE, 16'h00FA, 16'h000D,
 16'hFFED, 16'h001A, 16'hFFDF, 16'h0027,
 16'hFFD3, 16'h0033, 16'hFFC8, 16'h003D,
 16'hFFBD, 16'h0148, 16'hFCB5, 16'hFD4E,
 16'hFCB0, 16'hF450, 16'hF2B1, 16'hF44E,
 16'hF3B4, 16'hF74A, 16'h01B7, 16'h0048,
 16'hFFBA, 16'h0044, 16'hFFBE, 16'h0040,
 16'hFFC2, 16'h003B, 16'h00C9, 16'h0133,
 16'h00D0, 16'h002F, 16'hFFD0, 16'hFD32,
 16'hFCCC, 16'hFD35, 16'hF3CB, 16'hF736,
 16'hF3C8, 16'hF43A, 16'hF7C3, 16'hF441,
 16'hF7BC, 16'hF846, 16'hFFB8, 16'h014A,
 16'hFFB5, 16'h004B, 16'h00B5, 16'h014B,
 16'h01B6, 16'h0249, 16'h01B7, 16'h0149,
 16'hFFB9, 16'hFD44, 16'hFCBF, 16'hFD3E,
 16'hFCC5, 16'hFD39, 16'h01C9, 16'h0234,
 16'h01CF, 16'h052E, 16'h04D5, 16'h0129,
 16'h00D8, 16'h0128, 16'h00D6, 16'h002D,
 16'hFCD0, 16'hFD32, 16'hFCCC, 16'hFD37,
 16'hFAC6, 16'hF83D, 16'hF6BF, 16'hF745,
 16'hF3B8, 16'hF34B, 16'hF3B3, 16'hF14F,
 16'hF3B0, 16'hF450, 16'hFAB0, 16'hFD50,
 16'h00B1, 16'h014D, 16'hFFB7, 16'h0042,
 16'h00C7, 16'h022F, 16'h01DC, 16'h0219,
 16'h00F1, 16'h0005, 16'h0006, 16'hFCEF,
 16'hFD1D, 16'hFCD6, 16'hFB36, 16'hFFBF,
 16'hF84B, 16'hF6AC, 16'hFB5D, 16'hF69A,
 16'hFB6D, 16'h008D, 16'h0078, 16'hFF84,
 16'h0080, 16'h007C, 16'hFD87, 16'h0077,
 16'hFD8A, 16'hFC77, 16'hFD87, 16'hFA7B,
 16'hF883, 16'hF780, 16'hF77D, 16'hF685,
 16'hF879, 16'hF789, 16'hF876, 16'hF78B,
 16'hF473, 16'hF68E, 16'hF872, 16'hFF8D,
 16'h0175, 16'hFF89, 16'h0079, 16'hFF84,
 16'h017F, 16'h017E, 16'h0285, 16'h0478,
 16'h058B, 16'h0672, 16'h0591, 16'h046C,
 16'h0596, 16'h0469, 16'h0597, 16'h046A,
 16'h0094, 16'h006E, 16'hFD90, 16'hFA72,
 16'hFD8C, 16'hFC77, 16'hF785, 16'hFC7E,
 16'hF880, 16'hFC82, 16'h007C, 16'hFF86,
 16'h0077, 16'hFF8C, 16'hFB72, 16'hFA90,
 16'h006D, 16'hFA96, 16'hF868, 16'hF699,
 16'hF767, 16'hF398, 16'hF36A, 16'hF295,
 16'hF76B, 16'hFA95, 16'hF86B, 16'h0194,
 16'h006E, 16'hFF90, 16'h0172, 16'h008D,
 16'hFD73, 16'h008D, 16'hFD73, 16'hFC8E,
 16'hFD71, 16'hFC90, 16'hFB6E, 16'hF794,
 16'hF86A, 16'hF799, 16'hF763, 16'hF3A1,
 16'hF35A, 16'hF2AB, 16'hF451, 16'hF6B3,
 16'hFB48, 16'hFCBD, 16'hFB3E, 16'h00C8,
 16'h0032, 16'hFFD3, 16'h0128, 16'h01DD,
 16'h021E, 16'h01E7, 16'h0114, 16'h00F1,
 16'h010A, 16'h00FB, 16'h0100, 16'h0104,
 16'h00F8, 16'h000D, 16'hFCEE, 16'hF816,
 16'hF7E5, 16'hF720, 16'hF6DD, 16'hFB25,
 16'h00D8, 16'h002B, 16'hFFD3, 16'h0030,
 16'h00CD, 16'h0135, 16'hFCC9, 16'hFD38,
 16'hFCC9, 16'hFD37, 16'hFCC8, 16'hFD38,
 16'hFCC8, 16'hFD38, 16'hFCCA, 16'hFD33,
 16'h00D0, 16'hFD2D, 16'hFCD7, 16'hFD26,
 16'hFCDC, 16'hFD22, 16'hFCE1, 16'hFD1B,
 16'h00E9, 16'hFD14, 16'hFCEF, 16'h010F,
 16'h01F2, 16'h020D, 16'hFCF4, 16'hFD0C,
 16'hFCF4, 16'hFD0C, 16'hFCF4, 16'hFD0D,
 16'hFCF2, 16'h010E, 16'h01F2, 16'h000E,
 16'h01F3, 16'h000C, 16'hFCF4, 16'hFD0C,
 16'hFCF5, 16'hFD09, 16'hFCFA, 16'hFD01,
 16'hFD05, 16'hFCF5, 16'h0011, 16'hFFE8,
 16'h011F, 16'h01DA, 16'h022E, 16'h01C9,
 16'h0140, 16'hFFB6, 16'hFD55, 16'hFCA1,
 16'hFD68, 16'hFA8F, 16'hF879, 16'hF681,
 16'hF784, 16'hFA78, 16'hF78A, 16'hFA76,
 16'hFD89, 16'h007A, 16'h0080, 16'hFF87,
 16'h0071, 16'hFA99, 16'hF85C, 16'hFCB0,
 16'hF842, 16'hF7CC, 16'hFD27, 16'hFFE6,
 16'h000D, 16'hFFFF, 16'hFFF5, 16'h0017,
 16'hFFDD, 16'h002D, 16'hFFCB, 16'hFB3C,
 16'hFABE, 16'hF846, 16'hF6B7, 16'hF74B,
 16'hFAB7, 16'hFD44, 16'hFCC3, 16'hFD34,
 16'hFFD7, 16'h001F, 16'hFFEB, 16'h000A,
 16'h0100, 16'h01F7, 16'h0013, 16'hFFE3,
 16'h0226, 16'hFFD1, 16'h0038, 16'h01C0,
 16'hFB47, 16'hFCB3, 16'hFD51, 16'hFAAE,
 16'hF851, 16'hF7B0, 16'hF74F, 16'hFAB3,
 16'hFD4B, 16'hFCB8, 16'hFD42, 16'hFFC5,
 16'h0034, 16'hFFD4, 16'h0025, 16'hFFE1,
 16'h0017, 16'hFFF2, 16'h0005, 16'hFD04,
 16'h00F4, 16'h0112, 16'h01E9, 16'h021B,
 16'h00E1, 16'h0122, 16'h00DC, 16'h0127,
 16'h00D5, 16'h012F, 16'h00CD, 16'h0137,
 16'h00C6, 16'h013D, 16'h00C0, 16'h0043,
 16'hFCBA, 16'hFD49, 16'hFAB4, 16'hF850,
 16'hFCAC, 16'hF858, 16'hF7A3, 16'hFD62,
 16'hFF99, 16'h006D, 16'hFF8D, 16'h0078,
 16'hFF84, 16'h007F, 16'hFF7F, 16'h0083,
 16'hFF7B, 16'hFB86, 16'hFA7B, 16'hF883,
 16'hFC80, 16'hF87D, 16'hFC86, 16'h0076,
 16'hFF8F, 16'h006B, 16'hFF9C, 16'h005D,
 16'hFAAA, 16'hF84F, 16'hFCB8, 16'hFD40,
 16'hFCC9, 16'h002E, 16'hFFDB, 16'h001D,
 16'hFFE9, 16'h0012, 16'hFFF2, 16'hFB0B,
 16'hF7F8, 16'hF705, 16'hF6FE, 16'hFAFE,
 16'hF706, 16'hF7F8, 16'hFB09, 16'hFAF6,
 16'h010A, 16'hFFF7, 16'h0009, 16'h00F7,
 16'h0208, 16'h01F9, 16'h0205, 16'h00FF,
 16'h00FD, 16'h0107, 16'hFFF6, 16'h000B,
 16'hFCF4, 16'hFD0E, 16'hFCF0, 16'hFD12,
 16'hFCEC, 16'hFD16, 16'hFCE8, 16'hFD1B,
 16'hFFE1, 16'h0023, 16'hFFD9, 16'h002B,
 16'hFFD2, 16'h0031, 16'hFFCD, 16'h0034,
 16'hFFCA, 16'hFB38, 16'hF7C7, 16'hF83A,
 16'hFCC6, 16'h0038, 16'hFFCA, 16'h0034,
 16'hFFCF, 16'h002D, 16'hFFD8, 16'hFB22,
 16'hFAE6, 16'h0011, 16'hFFF8, 16'hFFFF,
 16'h000A, 16'hFFED, 16'h001D, 16'hFFD8,
 16'h0034, 16'hFCBF, 16'hFD4D, 16'hFCA9,
 16'hFD61, 16'hFC95, 16'hFD74, 16'h0084,
 16'hFD84, 16'hFC75, 16'hFD90, 16'hFC6D,
 16'hFD94, 16'hFA6C, 16'hF893, 16'hFC6F,
 16'hF88D, 16'hFC78, 16'h0082, 16'hFF86,
 16'h0071, 16'h0098, 16'hFD5E, 16'h00AE,
 16'h0246, 16'hFFC7, 16'h0227


};

logic [17:0] player_depth;
logic player_repeats;
assign player_depth = 18'd8731; // same as numbers of samples
assign player_repeats = 1;
/* end player explosion 441 hz*/

assign dout[15:0] = player_ROM[adress][15:0];//16'h0; // take the adress row
assign repeats = player_repeats;
assign depth = player_depth;
endmodule 