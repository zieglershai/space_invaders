// System-Verilog 'written by Alex Grinshpun May 2018
// New bitmap dudy February 2021
// (c) Technion IIT, Department of Electrical Engineering 2021 



module	bonusShipBitMap	(	
					input	logic	clk,
					input	logic	resetN,
					input logic	[10:0] offsetX,// offset from top left  position 
					input logic	[10:0] offsetY,
					input	logic	InsideRectangle, //input that the pixel is within a bracket 
					input logic playGame,

					output	logic	drawingRequest, //output that the pixel should be dispalyed 
					output	logic	[7:0] RGBout  //rgb value from the bitmap 
 ) ;


 
 
localparam logic [7:0] COLOR_ENCODING = 8'he0 ;// RGB value in the bitmap representing the BITMAP coolor
localparam logic [7:0] TRANSPARENT_ENCODING = 8'h00 ;// RGB value in the bitmap representing a transparent pixel  
logic[0:31][0:63] object_colors = {
	64'b1111111111111111111100000000000000000000000011111111111111111111,
	64'b1111111111111111111100000000000000000000000011111111111111111111,
	64'b1111111111111111111100000000000000000000000011111111111111111111,
	64'b1111111111111111111100000000000000000000000011111111111111111111,
	64'b1111111111110000000000000000000000000000000000000000111111111111,
	64'b1111111111110000000000000000000000000000000000000000111111111111,
	64'b1111111111110000000000000000000000000000000000000000111111111111,
	64'b1111111111110000000000000000000000000000000000000000111111111111,
	64'b1111111111110000000000000000000000000000000000000000111111111111,
	64'b1111111100000000000000000000000000000000000000000000000011111111,
	64'b1111111100000000000000000000000000000000000000000000000011111111,
	64'b1111111100000000000000000000000000000000000000000000000011111111,
	64'b1111111100000000000000000000000000000000000000000000000011111111,
	64'b1111000000000000000000000000000000000000000000000000000000001111,
	64'b1111000000001111000000001111000000001111000000001111000000001111,
	64'b1111000000001111000000001111000000001111000000001111000000001111,
	64'b1111000000001111000000001111000000001111000000001111000000001111,
	64'b1111000000001111000000001111000000001111000000001111000000001111,
	64'b0000000000000000000000000000000000000000000000000000000000000000,
	64'b0000000000000000000000000000000000000000000000000000000000000000,
	64'b0000000000000000000000000000000000000000000000000000000000000000,
	64'b0000000000000000000000000000000000000000000000000000000000000000,
	64'b0000000000000000000000000000000000000000000000000000000000000000,
	64'b1111111100000000000011111111000000001111111100000000000011111111,
	64'b1111111100000000000011111111000000001111111100000000000011111111,
	64'b1111111100000000000011111111000000001111111100000000000011111111,
	64'b1111111100000000000011111111000000001111111100000000000011111111,
	64'b1111111111110000111111111111111111111111111111110000111111111111,
	64'b1111111111110000111111111111111111111111111111110000111111111111,
	64'b1111111111110000111111111111111111111111111111110000111111111111,
	64'b1111111111110000111111111111111111111111111111110000111111111111,
	64'b1111111111110000111111111111111111111111111111110000111111111111};

 
 
//////////--------------------------------------------------------------------------------------------------------------= 
//hit bit map has one bit per edge:  hit_colors[3:0] =   {Left, Top, Right, Bottom}	 
//there is one bit per edge, in the corner two bits are set  

 // pipeline (ff) to get the pixel color from the array 	 
//////////--------------------------------------------------------------------------------------------------------------= 
always_ff@(posedge clk or negedge resetN or negedge playGame) 
begin 
	if(!resetN || !playGame) begin 
		RGBout <=	8'h00; 
	end 
	else begin 
		RGBout <= TRANSPARENT_ENCODING ; // default  
 
		if (InsideRectangle == 1'b1 ) 
		begin // inside an external bracket  
			RGBout <= (object_colors[offsetY][offsetX] ==  0 ) ? COLOR_ENCODING  : TRANSPARENT_ENCODING; 
		end  	 
		 
	end 
end 
 
//////////--------------------------------------------------------------------------------------------------------------= 
// decide if to draw the pixel or not 
assign drawingRequest = (RGBout != TRANSPARENT_ENCODING ) ? 1'b1 : 1'b0 ; // get optional transparent command from the bitmpap   
 
endmodule 
